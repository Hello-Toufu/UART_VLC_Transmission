��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)ND��0Ps��� Q�:�!�2�q����u0P�(ng�z�B�q�c�ld�lf��t��L��8�n)j�wVl�	�n�Ϟ5G7)O��_�ۘ�a�[4����@, x5k��(S����[��,e����y�����6�r<��D���ߴ�-�v��5앐4&���P����V��	�PC����n�b��K�GS��,��j�d�2���ث��?�&#Y����6����* l�C�3;ډ��p��;�找�ey�Ӡ���~�zz�j��`��Az�_.�����)�&�d����7h����)U�
JR�>jӍ�̴۠mB�����`��ք�;w�����V671}�|����$Ļ8X2qd�%��]ǰ�\z�^��	i�P�ۙX¢��N�
��)�{��Y�g�~J���p�yV�9�9��w���)m��_�*s�|O��
y+���MhF�]Ƥ��#=<��(�T��2�a8v��S<�}�?7�!��Z�����L�g�*h��}P'�	Eމ,C{�CQƑ.�'��a��c[d���h���8ڜޑ6`i�K#��}���3�jM��v�3-���O�Nq�q4�zJ։��4�^�o�P��c��v�.H���Uv�g�w�'� �E6�6�E|f{��ρt�#���`�N��s�pqSա�u<PE6��FgK�7@ڛ�Qk����ẏ�����F8�*�c1��3�3�N)�8Xbj˒=:g��Fo�2�d+�2;�i UK�_շ+o�s`���D��K�m�/����Эk��7 [����y`ߩZ^9L!���ά���~�K��Lˉt�hd	��ΌQ��6�X�i�CGhX���r����Di4~ofi]ƃو��2�o��4C��	lp������8��Q�d�'�Ӄ����{9�A�n~T�~���wd�C�u�k�gԓ&6Uyi�-�Vg2T�軃�� ����̳����E�x��4q���*X�Oy�Qi9S�bE�kqmc.yX��r��#����V�����+ ��5n5t%9�������������'| o���Ti�i�O��ma����\��xY�4Bwf��2��,e�$	<B\_�y  ��g��ZD�_�(�Q�MٲH%�%L�	3�໔o��;-�1�D�_Z<�����B��k��Xz��9�����ϕ�����3*�>A��?{��?b�fy�Sd/'0C6=<}L�(��\����0Q��?C�ط��� ���j���t?7��Y�U�