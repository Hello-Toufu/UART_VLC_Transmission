��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��P��=:� ����(�)3�� 5����l]0�ك[�Y�qޡ�(���fZ��#b�}a�3�
>cO��o�LW��4�C���(C��&{��"�v11#/I�&�)�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_��r��)����%|j��)����kMd{'��_�$�iC���ff܀���o��|��y�Zt7�ׄ�'抰�i�o"���MQi�n$�w�3,�
�r�%l P��l|�M�0a�ha��n������|��!<q�Ф���QG�M���ȝh��t�)�����������=�J>��(�4�b�^��IN���D0t���1-Z6M�
�*s�2�v��/�p�����Z��ý�����C��.�:��h]���>h&5�e�������t�;2��_���s���H�F���j����6B�>;'��g�z^1sLn�IzSg��en�?�k :�,�T��<B��T^�����s=�,lqbE6��*ޭh�u��p?�>���.ՒG%��h>�x��<�b�j:��/�|E�@9�Z�jk��I����8�|A�Ļ:j)��]�R���$!@�Är��zN@��C�Q�n���6��������9�_AZ*���Q��o��b�S��y�ⶍ��%������kE�C����𔭜!@A��Huv���2��CĒq�V�`ͣ�stY_��^Q$�y}<�X����
�%���:b�~+��Z��h�N��/��+	���^��4�&苇�]�~��W������x�y\��%>��c��=��+���9��_Q��B�n�}]��J|����ʿK~U�i��%�X�S�TJ�"5�_�M7k)5��ZN{;O��������@�YB�����������ɖ���!��n�tI��P��x*��&�x�?��Ps�9�������9'XX��؟����NCF�o�R#����x��_	Ѳ�F�