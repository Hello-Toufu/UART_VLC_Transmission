��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��P��=:� ����(�)3�� 5����l]0�ك[�Y�qޡ�(���fZ��#b�}a�3�
>cO��o�LW��4�C���(C��&{��"�v11#/I�&�)�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_��r��)����%|j��)����kMd{'��_�$�iC���ff܀���o��|��y�Zt7�ׄ�'抰�i�o"���MQi�n$�w�3,�
�r�%l P��l|�M�0a�ha��n������|��!<q�Ф���QG�M���ȝh��t�)�����������=�J>��(�4�b�^��IN���D0t���1-Z6M�
�*s�2�v��/�p�����Z��ý�����C��.�:��h]���>h&5�e�������t�;2��_���s���H�F���j����6B�>;'��g�z^1sLn�IzSg��en�?�k :�,�T��<B��T^�����s=�,lqbE6��*ޭh�u��p?�>���.ՒG%��h>�x��<�b�j:��/�|E�@9�Z�jk��I����8�|A�Ļ:j)��]�R���$!@�Är��zN@��C�Q�n���6��������9�_AZ*���Q��o��b�S��y�ⶍ��%������kE�C����𔭜!@A��Huv���2��CĒq�V�`ͣ�stY_��^Q$���j/���I�N��[�¢
��.�Iǋ2�RW�1�X3N�~��p6˰b���.�aS�і2`�C�	o�߮��ˮ7�/�ఔvŁ��PA�	��>���>��f�lr9T� �������t���Q���;;���*A�0
�.��q��C���*i�ZM��k6|T�&!��Y\V2,����17hsE@���:�k&��CR@ذ�k3�mqM\��P�`�FӖK�V֡fˉ3)��N���$'�ԿW��q|�8���Ĵ�'�E��Y�T湥��7zr�e��K?Ƽ�c�}�b��F�G
 �z�"�7����=.�~.}��B��H�	s��\���}u�L���.��"�9٬-�m�J9:��:�:	}�:��R��L{a�� 
��Sʍ���* ����`��G��9J_��f�j�f������<�~2����`�,TbtBž�A�����ڏ������ -����r�oz�6Q�{�c�]S��*�n�ָu��#B7t��u��좠��/i�|�W7J�_�e�1���Fq:*�A���Ų�]�pG�ْ8oQ���y�r�͌���
 yW�R�ɸ���fA��F��JC�4޻���~��@rA~���nO(Л�m�}�cI&�!K�¾n6y��݁��[�A�\��lv��:9������<�r��Z5��W�̶<[9�)	���@�"��w�a��$��Qm��QIn�����Q-�b��/�Σ	җ���-m�*� �>�D�M�o����|' ��<��*��y�.�Ku/s��pfX``��q`�]��z|R�B-����f>y��`��z�ؕ�'1�Ba�mWyX��b�ḓ-8�N#���Y�=~@/t3ף
������Lڡ�v*<R�[����2M�m�|L�)���:���E&N|zƬCe$��(�Rnm���$�)�:5�;��q8Jd���C��ߵ�6��]��I�<�-POƴV�]�R$~�GY���i �c��f���`W����SSY���h�!&��ޙ6��3���j��p��|��HOBG9>��_�r�@�0cP93�F�*D��2$U/F ��|�h6�!n�R7`�;�蚬v��)��l/Ɇ���%I�g-й�L��%�l�*b[bE
�^�@�c���%��c��BYyk��y�/y�� d�z�����eO���)=�0[��d�2S��~j��,�}<�U�"�p	j͊�C��Z(#1���4*�J�,}���������<��W��h��&��W�2QԻG� |��J/5��Ѯ�g�Tں�G��E+�!�3�m=�k3SM{�d�4EHƟ���?a�R#,@7��Zl�h�`D��aGS����a�{%��ź5�	*�OWHl���X%Z���3xm�xSҾ{��&��@<\