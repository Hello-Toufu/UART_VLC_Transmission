��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N'�|Z_&i��N��wG�����=p�v\G�;����?�T �?þfᚶ��- �r��6�mro)����'M~T'�6k@3?�5l�&�\�< :�ڱCs���-�5��-^��6i��S~���'Q�!ݫ@]Q�Lu\u�G��u� G: ��19�selG���2�J���B�M컉�s;܌f!�U?䥜�}���xV�������h���@���(��Ys�%�k*��$f�`��9��|��Y�_�.��x�Xf�@�U�j\R�H�9�����-PlA��9{LMR��Z]O�ڨ;[B��|_���8�aZ5�g���i_����躆�����SL�h�7ï��ݰ�k�����U��ԣ��.͐��o��}#�0��}���	J��3	������7�J��o6p<:Z#%-8+��w��3T��g5��y���  �����>Evm��w,&_���z�e*�1�-����][6�q�������`M�Yq��!9Tf�&��/|4�)&���g��;BIA���lʘ�4c�(b�`W�2�;�[�Պ ��z�S��nؔ.��M�}'_V79���ϕ�}�1LK䐚�s��Ga��sAZ������Ū�;<\o�EavQ㸕��5�8��=	���2�[���hD}�!Ԅ*C�Iy
��%4b�].Qi��*1�wF<訶#1i2sZ;`	����u9�r��} �p����n�D���@��lw�ǆ^�6�MI�[�`��
*@��>�,�����~_��E��N;2f��d�j-K]���Jj���r�#ꖶ���c�??ھ�IhQ;Ņ3�*'�x��{x8�]�ٌR2�-��=LD�}_1ظ�&^*d��K[�'-��!�����d�_�q+��YP��ʲ�	qpǑ�P=��=1�`\���o�3���:���UyNxIV�S�TD � 
{(+�#������!Qb2�������ӅI
t�����S�0R�� d��o�KAj����`�p�@Uշ��~#�;3����;�6m�}��3�^M�s�2����C��9� �����Sd}I�H�$�}�LHʰn@�j]8�F�t�������7���o��Y�(��Ey�_��?���"�H'���J?��e� _P�	7J���Z��^�%7�a�^���l�H��V�qv�L����䘔����y�A7{�X��7�Ԛd�|Y�P�4�c��[Ȯ����ݡW+�/S��8wF���s�~(��5d#�m��$�i��7K�}�z�G^C&��