��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�G��ˊ�I�2�8�D�ĉ�a��{����[�^�ڝ��m!��
0�mt��|Ew@6 0(�:�L8���A'fܴ|�!p�詝�������~b���&��bL� �oR4���U%Ы^��<�dC������+�I媭�'fB���7LO~k�
��t3���be���t7a�3��z_�ܲ6�~�U�JaQ*8[��1�Y��̬A(=�D���M|�^
���M?�I{�/���6���� ����h��I=�O�'���4��j�gʳ�X�+�� �1;�8�ݶ�	n�X�L�4h�[��}���M榞"�IS�7N~��Pkg%��I1��{�����a5������E��p|>���<+Ӝ؁�5��؟.A��xE����+�0/�����OXBn���%D�Fj�c�h��7�W����>�ͮu��]T�>Z0S�n2�N0>���U�EBpbWqxg"~:&u�0��`Q���܃���Ǒw-��M���D����u�\����g'���E,���å �J�8F``��	�C�����6�����bi�_�J�����P�ʐ?y� J��ٕ-�$ 1z=�If/� ����3TQ���+b)�1����I�����j��YLm�HKT�N�����A��(ӈ硊QI6��3���M��S�����m�aZ�'����9ą�u�ᅸ��1♻)`[�V{��� -��%[��� -�unG���8���&�a7��kW�=�:6�l���6�$�o���Nᰱ
��L�M��M�$�!In����yӫk��*�(�&�<����7X�̩Iӝ+ �tǜ���k�hIm8Y�C����t~c3G���r08@&j���}~D�ہ8�B#��`���Q��9+`/̩?�ls{y��'2��MCWk�M�\��z�axe�O��C�H��)��`�7��=i��