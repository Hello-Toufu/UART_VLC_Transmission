��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_��Ջ
i�xH�	��P�������շ��.R�a�}�S�C�+2f��l��@�I �1D���9���Òz
�G���` �㑅sy���C�M��"��	Pp�?��GSS
2$ŧ:F������'z8��ѓ�:La�olFZ=��'L�oc��x�!U;oܶ�xd��G�D]V��"B��d�m�Z���e��{�����]'4��۞R�_-ʗ�T~��y�RL(�g2��?�j����Oj�4s9 Xv��t�� �IEn3S��Gd⬾
�5�p�+JQ#�f�0��YQ�8��//0���p�\F_�wimMcl�=��t���>53���]�hdz.��
<k��t��8É�|8psW��mszI��D޿e^Oo��t�Q�|���)Z�c����C�[����ͯK%a��3�G����KR嗬El�`b�l�*�O	X��)�J׉BĠ��l��h�1�R2,�D�x�bWb�u��rl�s��:�K�)իp^�O2�N���A�(����/���_�Б��x�.ld�$�����it�J�e�*%z�!�+��&�AJ������@�9�)=�
A�~\v�Ld�\:/9W�U.w�B�i� Ŗ�hr��(�K��7,ye��h�F���	6~���u�w���ֹW?�J���:�� ����k�5(��s�͕|N����v�,���3���EAD�/����9^�.OZY�-�D@Ķƭk��6�Jy&'<$a���@$:�d'30�P��0�K�rH�*�i�f������O��_1�_q�ܩ����(��������ql*��!x	Q:��W[�|L<��u�����V��`�xW� +�� �\����oڱ����Qi���pT�{�bH�w*�`��{8�U 2߄��_ �E����ZaN�m߼^���[���-gL��S�-6�Ď&FM$%��J�'�@�җ�։[FF@���1�3'1 ��*-��)��)vz�U�">�zF7�\ �jr�2-sᓙ�)�^�:��3���CĤ��淴���w�����B�pl�w��t-�?��0��'��U՚�z9�W�����|?�X#��5�ܦ9�ו��z_�?���cFΠ/����3d�D���w��ë�o+H�_����m�=����uK���N�!�BY���OH�Q�#�E����MA�jK��q�7�M��M_�t{@���)l�����fQW� �M���@ ���E5��;�d(��.���ֶ�0tk: ���#��gz=+�����a����l��R��Y��m�9��"�{T��Sz���<�˻8�;Ë��Ә�a�Ƥ:_ѧxf����H���o$���	�h�ٛ�=���&�T,�䢦+�g^ג�1,3����?��3�a/��>*?����3���=&����.hRu�e浫�y�Z?�\b=�{��\��Ah��D[�Hjl��n�W���yz��`$�(��Ҧ�<�W�#?x(�M�������s--�ޭ��Mu�4.�k��q�8o:䃋��c����kSg'�:-<��ˊ����5^�7
l�s��9&EA#��c:���R�c��Mެ�S�f?��^# �2}�����5"a�}ӫt~[6|�0�喙�'3#�H��Ӹ~1tN�BLz�
�^Ĳ�l�M��+�ƙ�i�k�/xs�C ęH�q)�A ��*VN6�Y�r�/p���>�{��� &g�ʅ��єbsB�9�:�p�y%-N\H6�R5�F�,!	���lS�����7$k�C�u����qL�}2�`�L�VnM	bp��S�w�D.ޝ�P�{�%����*a�N�v��8�����5c㰗u-c�dR�:AQ�s|�!�dZ �-ke2�o�P��=Zj�9���V��� ��Ag$��w���DFL���p��7����E�/"�X��eR�w'��$йg���;�q�'��"�L�z�����e,�Τd��=�+!�hŲ�L'����d_=����hg�>��\����@�����e��ղ�Z���I�*��d�`;:� ,��d*?zG"����xI��h�(��c�`ѝ%��ʂV�V��3��ݜ�-&����,O������P}*a�:8��mT`����@�7kj���Gj�c�)0��z�����
��pa!�#8����<<x��=Z���Q��^켚�����֢��II�r��m��Z-�y��N\����k�UqkX)���>�B�^�pc��^49�����Ca3�n�S��s����N�2�i�R�`]�˜�y���`��\�,��ܒ��`�9�S����$�~���rU������A��ʽYց6t��o��r#�'��އ�<#�=��9j�"��<���I��#5����
�kԓE��_���i "E����������Fp�a��� �jC	Zƈ��yo������f�:�Ԅ���wu�BG�]���9�
B'�3���Ũ����|[�&AO�A �\�!1;��𗁆�E�b�T�R�
�AJ�wR��}+���� ��"-fO!B�C,�s����Eۯ�2��kt�94Q�B��%V(�p�D�am��l�TB���⼥I	��?o}a{\�4|s|?�.tX�ցZɥ_c�����XVcSir�gw�}��
��E��gS�N���V�ŔiE]Ũ�X-��F��6˱��Ce/+�a؁�K�LKΓ^�֬�6da��A=LL�U�ɏh|���Y�{Y����p
���`����H�=��p`�Z{H���8M$�:��?�Mc,_t>"Ԃ�Z��`��'2�pc|�w.c�V�j՛����A!�p���^cJ�?�M��YN�����,;w�-{d�G��K$K��*��3U�)�:<�=����8O�y�F�(�Z��4�qx@u7jz{��J3����̤�UY�.���S�����
-�᪫�U�d���~؅^�f��q,��}�8
��qΝ%]�0�W7��ኳ�ʬ�~���	����gdC��Kp���f��fe��!6R��d��;�VC��C�kR��y���*w��VQGU�e��F!������P������$����Yx���$F�NPf�gɽ��C�&�:S��B\�0%@��࿬a�<�3�۳��<��g���W5-�:����2��~�)���R�%r�<���c�K�0O�Au�k�l�KUT@���%�����b*������!�ZPW9S�V[�������X���p5�7��+R�XT��&$���~�0�����ecd�,;sZ�߆�)��0 �����C���f��gj�۴�D�׾��so����K��Nc��I����'mJoC��m!��6�r*�ĸE�Vz��R���*9�7��c�m���,�n�a ~�4+��Uc�������֝��W��F����O$̝���(��`�8mtمKiS3�ٝ����Q�	s垎�L�Q�����9�k�s�8�vx�(f�r[��KT!0a�S12��V�� �)0�H@��DF�1}Rvw�1t���G-Z�IMpgL�G��Z��2`_P5��Ļ�C�r��z�7v�,��y�{�}Rz��ϗ��gڪ+��ǫqҬ݈Y���Bb*Ԩ� �^.6 �W�)<����=p�1&7��׹I��p	��b���X�(؏��H�uؠ	��g�	��V���~��$��8h���w�X�S"�d`7z�:7�j��6{�3�mL8Ű)��p	��6���l�\ä7�è�: Ĺz��-"�u1�M���ev�NbG�1Y���z:|�fg��ĈC|��a�S�OJx������:�M���A�g�&�VI���Wќ�
��O�㡒sХT�"ID���M�G�pڷU�]au(a�Ɔ�d��.��H3��T?�%�9>L\� ^���wR��;��!QIA�9�ŧEcc�ןN��aC(A�ª��`N��5��{(j���W��MZ�A��V�s^���S�2�����=mo!�Rp@����������'���P��vp$�T����x�y���8�IG>�h6�o"�
���=�ޑ
�h�"F(��� (�Ҟ�)_���8�F�6��dB���3����	�l��J�s�\ث`3����c��Tl���ރcɉ\jm�ˈ0(�\a�k����o���@|y$�r��
��n(�|:�����$��<h���"�d��_��$ʞ�IhXMEh��S�	Z6x�/�X�z�Ͳ;0�x
��p�$s%Bn��k#��=�E��N`����o-��
�u <O0�k�+%;l_}�-w�qx�������g��=
�>���[��60�K����ׁ�����,�w<w^[i�h�7����+�`0�3�.��h���0��Uu#�O�����x�alx[�+ݷ�����r�#�_�n'���܁9#���F��.�t%s8z��	����q�*�Ρ�+{ıw�T�7bUBdCP�jX���ެ_	Z���8'�s�$ُ��O���=E]�@qV�ބ8���,�B^s�ͯ�孴�a�~���&9���|��5���t��1(���3=�A�T=R<���MY���\��%���p
�k�G5���.r�	^crB���qM����n%خ��sҝ���#�lQĞ�[h�c�[�@~+Շx���� �@�L;lgw=���B�w���F����D������!�$�l ��2�b�<��)S.�����m��WǮ
�>�����V[)�e"�Dă<��s?��&�� `x-���ї��2u��rq��n���U����z&��X��ǁ���fxޔDM�⡸�����{��ۋ�◽�aE�S�"f�^Zc�J��9�a*������*�B^��(=I��ڟ��_��3�Pf\_���68�'��̙�k{]�e$���e~�nk[�w
��H�G{0)]���h���|�.�t��"	�T�԰5K6�8���H'��tPZ��-<yc�<��׉m�y�j8?	Pݘ$���\���>)��;G��C��`��������Q�`�@�W���0}�b�4X�H'Y?��[�S��e��5;��=�p>>���`�]���\��]B�Vt@#�E��&��h�1c�6s{��*�O-!��6D�B����)�޵����$�v�D�6�c�P��Δn"rS�<OL���M��@�����4���vD���^D�ܺ�؏7e/J��Έ�ɒ��}H���{�D��B� ����(�M��U�+��q��L��}��I,N������帟���/�g~��<'0�pE�g�]�����Ҋ�)�ut[����>���m565��
��t�K�uˠl�6��^��S��?+�1�Ơ�2:W���~a����od����ۻê;�K��L"���V`����v�Ţ$&�[�1%)���0�)Pq�];*Ǚm�f`#��|�b)�k���c�K����IoI�247��Ow|��~k�<DC)n��e,]Dw)
h�_R�^O��+�p0���4#U�切yа���x2�NS�s(+R�o���[�.�r�p���R�Fd*��!�1Y���#z)��T� ���c�ѝ�E��H�Vɬ�i�,e@�I�^�呌�ǟ���c?��Sc<n4���e4r��<?9��AFdl�<0�k��Zmѽ�gO�~/(s8��n��b*���`��HRm]�e#���E8�����T�
9b铛�,w1e�W? 
�4܊'SeuN�*g=�����D�՞���'9�ƊkB�9MFc�Fݺ�ǰ4�&��R�����#*�60���&�vV����{����߷����c�О�FngD�#���ήH�M-�CBL�fB5�4K�2�x��
p*V��U���2�g�ng���2���=	N��%��������M��^���p����a��s��_�T:~�����Y����hy���I���D��&},~Թ��U�U -܀6�-�n�� �nX�#~=F��D�<y�"�����Vͭk��(��/��bas.�ZG�m=k�%��\���]8�ԞLz�:)����y�mŐ�%��r�Xt@�	��/�5e�b���;�����6Y�d$#�ШBz<
t�3���=�/8F�B|U���\��ك������7|�_ H�>CY%qq��6�����F�	���yua0��p�����/?�'�?_�jk���OmO�#�g턑z!�l��J>
��)9yV]�S��c�W����Sg��f�y' �Ԭ\$�2.���6����Tc�$&�jk��_;���^a�^_o�Y�_�{qT(�./�����֦��e];�d��.4��e�̏�w�{l���Y����H���q�mb���$,��5~6�*ƜCȏ�E�;Ƙ��阭�yT��/�r�(RR��[��g:��v���t�`�Z�&'��6�9��"^��k����+��Dn�t% �o��8?&A�Uv.HR��L��dÖ\o�D���g��L��|�l�@����c����u	�R���!khstEV�ި����z�@��ꌪ��u���O�e�P��aK��7�7�n ����_��x�/��(����#?�d��l��sf�.0y�T�O��5)�Of{���<ǦA�z����w�ʏq/kZ��%Z�{���r��ѧ��x�d���X�6tg��eC�Z9�sK!u��]C�݁nx˜���O���u/8�"G�I��\O�����6'
�8�c����M* ^����U��L�sX���(<�$B��܈�J␱T����6��4{җ?�v�ʕ]�V�,�|&ڕCW�1�����,
ji�D.ި�̄J�R���fW��fǩ�""$l�MRox�؀�y�>֌N�#��tt�:� ���DPh���S�`F35�窕�eD�?�G7�F�l��t��\{��2������8}�1ۨ�@�Ʒ.z�(4C_��Vo$�z��#�sx�?҂dx��T\�1E'|�i�`����A����i�����W�J��1��Aa'ռ���݄��W2�wPun��g�-B�/3���ӃkL��CK�W��и��6Gmh�NN���Ƴ�(�x�ԯ񕪴��#1�W5���S�N��|F�l����?���l�Be����-���&��������e�����7�׾�{ ��|�?�7z�ġdy'Ѽ1 ��*���\�2�ۍ��(|���:b��LxB���_��A�̇<��,��:���(	�Y�p�����q|������8^	�)�]꼕��](��G��h�P%h	E�w�B\z(����&�w��1��5;�� ���?��|��6#GkӗUK�U1�����0�rJ����(�G��j\���5;V��k��r��>�	�c�+�Ow�qj�z��Y2�O'	]�{&g4�2�J�T���߄Y���!��"��L�1����]��\��f�v�n~��!xG=O^��y8�zp�Ŗ��u��Ȕ�wh~5}�&�d���B���!��/Ʊ0g�J�$�b�cs��f���mz�����5���9����#&�IW�O�X����ȿ̲WT�ucn��,υ;�J*}�As1��9+}8Q�k���2��@w΄?�#.F��bow�-:����1��t�~�`��_@��M]2]��Dst��!����mHP�^���RW���
���V�!�W��\!H`E�h����ZV�9�Z��"s)gmwdx��+��v�Du�;C��F��������T�V��g��˶�?�����,��6��f�� ��i&�0i|�z�����͵�7 ��}�,t���\NSp��/�CT�5�{��gA��ƆQu�S��`V�
5R�/'1;��h�2����M� -������aѺ�����6�o���� 69Sz�O���!�T�͊8�#�ZU����WC�kv�w&��_�O8����6F�
�K	�2��Y����y��3�ZG��?o��OH���	���&�`���D�0?��[��Y	���7�Wk�,j�C���RO��PF"#e���.��C�1c�dj/��j��>�ly{��nD��eC['\�E�޵;)�j�Th�Ϯ_H���G����&B��S�y�·����o7cA[�D�j1��*�73 �p���Kب��xk;�1ؗ�)tJB���W��/7��`�R�v�J��fi�����������"��(S�k̑x���ރ�y,��ܞ����`��9am�%�J���e/��o�s�*�3��-~���L���@6*�R�<P�p�\�]W� �����~5
3�Q_STmسY�>E�@>a�?�J�t?kFj�bJS���PSu��2j�JG��
]_g�L�[>w�Z]�Y~HG�Mظ�C�x�1���bTE@�m5���6P�qF<�`4��k����	������z��W��U��_�,j}R�f�)k�%1�,��2Z	/�V�5�R����з�4u
*�X��K]CG�s���w�Y�z�c/j{�7'=�ed�ظ4��7!�8 }�j�z�y@�6}b2��+�(tiV~�
 W��䣛�{�{x�X�L��J�p�	�;���w9�{�#����@�a>�g�k�C�m�iDo���!ݵ�S,��+��d���{���O��
����䚮UA`2�?s5�n���U��#�]�Do$��/��t��f�M�]uKӴ�ƽ��ߐ�'��g��7��F�4����B�2� 9r�VB�zQ��rq��`�0��[�8Y��c���Ep`��(R�w�L���(CA�������o\�l�ޘ(n73h�$��JV���`{��k�U����e��D;�����F��3�qtPB=�'/�����iN�����X���G �s�evKrc�)��a<���ʶR�S �2	*P�DV�� j>���9���iз�8�j{V:�:�խ5���Ip��-_$�}��7v�:����Z��=c��~�����&RDӜ��.���2{<���w��bY��g���������J�t�>�A��?:2<>P��kk�_�
��;�\u�L����K'�!l�u�bF�6�l@ls�Ub�?�Y- �c��H�h���6"���� <Y.� �>p������h$.]�Q�iÓ� ;T��E#���/.���ﲜ3�:ol��xI�M'�z���#�O��1��5����7h-���їTc��+���x	���4�g�I^�#���şn��\U%�߼�pTz���`g~�Ww�> �`l~Cp��EOi���On}FUÀ�r���� �:C�ؚ�P��M��v���sB��gPFD���.�k踐���i�n0�Ѯ����g\�5��e��t	��~�:&�����?W�$�#�@'?�[#��	�3[�ԭ�T�ּ���=|� �̺G�U�Ȥn� ��.�X��F�2��=��wW�*q�O��Yh�Z��O����n��l�gz�f�*\kvgN�$�_q�I����
���\X^}���W���w�����Ь%f���`/�2?��j�����[n�'�u;�:�Է��Y��	]%U[n��m�I�\�˽S�����������g@��EHTUr��5�i 8���G/aJ�F�fR-�M�-���ۉZF�A3�����4��c�氁YK�0H��/n������ʻ��Ś#�c�[�8��j����Q$Y9̻�<�X!�5�:^��˧(�]mAf� ]�����Da%������6[�y�S
�G���Z�`}���r��+����픣�A��ʥe�Q͢����@�x��H��"z�φk�SVKS+�_���������P����ֽ�	�Lb���i�����
0C{�>�����!����ڷ�1��yi����2/R������aT�����OJ������(��]�����i.��0���Y՚/Ǭ`E���,�u�Mw��K�P�S��-���ru6]�a�@��Mr�풐���0m���`F�+��%�$��ʐ��g�Z��D����{�Z%�'��$+a/��؈�]�9�u�(�/ϗ_(��Qvb`<������Q]c�x��N	j���Q����������Kur2��O�����mZEe��w]R�9sU��_�)Ai��"d4A��@]�E�'�U�����k��\_����=�I�8G�z�s#�A�����!�j��0�*��g��v�f,�����K���Cϰ���ϵu�5� J[-li��&{�y�£���KDe]A�v��1[�I_��Z�|p��;wo��4#^.�xk�`�.p|���e>���[S�-,�Ȕ��y�N����	2$�&�U���Q�b~!$7�L�^s�NAQw/臆	D�2iY���5o��Nd�Պ��\�sNFSl(���Q�E��2n�������)�q���v�T�	7��D��t���QB�-}<�<B���Q
��f���hT�����4Z.b��U�Fe�0^D�	y±7J͗V�zN��"�\}m;^S���J����q�f�D�4_����ߥ.IJR�"�Z4�L��Q��#fwT��N�
���B��>���j�Ӄ��*��݈D�4�"P~u��qΰc3G��u؅�n���ʲ�C�;�9â�܉�],��@]r$J�����3�>d��v��B�%:I�5.c��Z
��z�_�!\pN㕾TTHl�) X���h~Y�=���gĜ����>B;�pم/%/m�	�9���B�������.�P[��əݶ�e����>��i��Գa���њ+�|����D�|M��
�g(�K��g���BD�q>� ?*��f|GKv�����x'����u�����y�sb!ҝ�c!X7�dȲ��;���L�I�a��X�� ȇ��Ȳ�禐�e,���� Z���^js4�d�X�#&aA�n���6Q����su�՛(�	&�{��9��AZ�𧉁��@u'd
�z^�cH�x�Vm�eR4v)�`�V�����/&ш�n�p"��x)y���%�^��z�18���#�O���u։�{�{�wi�EΫ1#	���,�VE�m�T�j��� ��DZ��رz���p��?��F������&ak�e��P �+���j��w��ɇ�a�gM���)���d;`�b�`�&(��'吋}�)���ً�]f�\9�yU�H9�z� �y����\�𐱙�	t�)r�*��ı9xL�bӸ�H����q���Ls��RF�-����o~���(Pk�W��,z��iO(�i�d��G�����E�H�k�a��e��Jt|�q��>�׵N�h�ߪ"z?7q<�-H_>/�����.����^fg	���wƜk�����@Cu��2�.{8�L͡�r�絉�rW,d`-�g�A�jُtEN��l̵�L w]�	��|f��Mq]wd���=�����/}=-ȧ����i�\)�� ��!��sNw�B�(�Ns�G!��g|��ak�ڨ�f������-�'��/QS��?�.#*�e�h�,�,Wr������P�X�j�"W���Q���M�h��pO@ 2�T Ï`�Ve�d��*3xA"َ7����J��k������F�uA�;�v$�7r����XEAv�wa�)u����_���P��&'uLh
�(U����H�ڦ+O]K���hMH����ֳܑ���'[Ā�vJ�޸��5 H�$o�HS���O��Q��V�gr/K����}�KA�6*oѵ�-<٥�pe��W�EoV�KE�Yk}�ld�}E��Y��a���&�������?Rbn5u�{rb��5�����&6x���0T�m3�jS��2G�tH*�'/i�*���&�����ܞ��[){�b��O�d�����I�B���өQ�A5�{�%��g�����
e��h�-O^�D�2��]ug<}c�fA�Ѻ-G��7.�e�S�2���[t<���ux;�e�S����M�U�R��y�m�s��^�'����5�E�sR*�#/jrˊ,�j�+*��p�����_YA4vGSJZLQ�(C�1�1Z�z���c~T.d��"�\1�{ѧ�X�:�9��6����(2,j�W�!TԾ�lvkn�~W��Q��9���%����u^��j� ��\�7~G���\
�GC�b�'9��qSR "��'�B�3��;JԀ��w䷵��	���+*(=&���/D9���J�3=!����3[�8��Ȥu�ڃ�����|�Xܑg�1O��7A�(w+hMͼ���`#�O1c��7�џ��$�ٌ��ы��)������n��ҼOi?\޷s�+���g�r3�k�s����(�M�|��^��t�vcڬ���lFn�o���i��
}�tb
~��LO | ��)u��*��ԁ���Si8t�Z?���2��b UA�2}�,�'�cg��nD8��$��Y��;{0�`?�ƝsE?ȡ26x�#�Ԗ��4:���V���曇ҿ��O�ER�4����&�����@��ƽ��m~f���R5^7ǝ�閡���R*f�R$��y�ױ���q傍��,n����� W���[s�+� ��=�C��5�I�n�2�L���a>���Q���Hlk��a�9�]���	#Ȁ	�T7�qN7��-��iG�׌�jݠ�E���H@�W;�>�	ye���(�c|���R�3K����o+�}���Gg�l4�4�7������I=f'�<��W�v���Eh�����'����	KԿ�S'>�Г�r�O�t����0�)��Ì�>d%�;+'*�b#��T��[��`�Gj�)���$#�E���Hx[����)���8xlMXv�޿F,J��W�M�ySͿ=��D5���W��Ϗ~�<���^|��O���=f0es��̳Lh���g۫T��2]w7����� MA�G (�-(�x��0Y��6�
0�.��a�Mu9�g�ӻV:�Z��%�B������\����+�6ԾD��yj�@�15}�I��6nᬅ4M�����<f�vm�.{��ZP���J�L&�Er��	-W��[}��؟�
� ��{��H,��$7̶D�C���p��|��f`�n`ޤj-��M2�}�t���%3�/1�0����8kq��z��9zn�T-���'�)ZԠ�+4�Ͽ���/����c39�i���C�0xgE
*g����!M��,dL=r�. ����ݣH���8h�V'�9?��P�Ԅ������AFY~��H1�C}f1ߟ�����3�fo�9�z��i��]���(����ۊ-"(��X��=}�_P͚"��e��W�+Q���-��u����\r���{�5�/�K��aߪ+1pg�o"D|Aj�����6��Y�s�/w�o��£ºs>U�N�1��a\r�k�΅�0�6es@Үn�XS�8�?�Qa8��=#ڌm��áڏ�b� u.zљDw���v�G�����rv;�	L���x"x���Q�9ǲ�0S���J�4�/'���\���dO���K�c����6�f�-�=�ס��𤋕T����﾿r��?S-%˽��:�Y�M`�4�֎�g�����K)I74ϲ'w#�I@��o"�Z����b:���#߼Vl�!]�s^z��Ӯ��߬�Ԡz����2��o��8 ��,Úw �Zb9A��G��r~��EoQl,�#-@��e��n,C��Z��P&��5QZn̒�����	�x�my�+nf�/����oM�)2v�GЌu,�$"���GP�}b����ݝ@N�|���x�X�r��pS�X�C�o�f�'��5���aP/z�4��}��/
e�1���*0)$8"hZAb�p�kTB�F�I�c!8��,�h�CS�F���;��m%�����Rƍno^�xO?����&D�;��~.>yJ}�u�l��|�e�H�A��G�nI�Ii�<���P��	�M��E���^�2�B%���1D�4�U�^�杩���ܖ���\��Ms��N6�8eRL�l��1���*
Tֲ��}μUm"	�`w�����Ti�x�p(��>�$X�F���(� B�lo8�N�����rK4���V;
�X��_χH�;+,%c�0X_�7�	vlf
��F�)�l%���D`����3���tG����^^ ���nE��C���G�գ�j�x�ϡ��鰊G�%��	߈�:`hiּz� eB͙��#�ބf��#�����Ϻ��Ȩ��+!�����E�+����<����P�l&�s�{f��F�(������Q��>r����+9�i��:��;�0{��>���}蝎�j��d��xȂ�콺�F��x
�5`�_3�}���h��Dd��%�y�Q r�A�(�3A_�2X�\�Xs+$|�Q���p�J��>���4�8+	8�.��DA
�>�lV����R��`�#J�Y�e��B)��|�E�vc �c����x3ة�eծ�,��ۘ�b���Q�h/Gs�%ǋ{��6U��!����K��A�(��%c$A
�q��b�U�Z���{<�q]�o�"Q�-Z�C�iE�!�˻p����7D�\y@Np�Z���\����r�* �tW0~� �Qku���`VA; a� ��Ơ�ՠ'�^�˱Y��0����?)��z@zۗw|=� ma��f��B����p|�by,���Ms M+<��FZ�xRF�TBCg^< �쯡�G�;BIA�V��w��.�]+(�t{��Ġ;��͟0��N��r���pA\S�� �fC�TQ��8l��	EgJgN��2�~YAx����!�~$�tt���p��u��	���hq���Mnc�^P|��d"$B�7�9��Q�{Ɨ/�:���qJg{9ͳ�0~���x4�(�+tnΆ�r<g��ŭ�Vt�=��UY�ŕ��7`p\��d���.oz�H��Ih��+	Z��$}����}��.E����]��6x�7���@�A���UH���<-��֋�7�jш���G@���{�=Vg=g[+^P��ϔ���&���.\0��!��P��Ϯ}�)텝�)y��B��ۜ�F�M�����)�սI�e�V~�h��SW�l�G�@��z�(���/:!
}����}6y�~:��D����@��E��M\K���1�ï��+��;� +�Rذ+wz�q�A�J���]�eU���p�^��:@�_�e����s��C��h��?꧟����zS�@�������P:�P��k\B���c��x�`Ds[ta?�?�Ȇ�{�r"����Q��wo>��Y��v*�����x4�O_��0�\��qZ�'��b��@%K1���p��C��VI�qSJ�Ʌ��a�h�R������*(�B�r��ţ5��N-���:�J�L7xc�c�ʒƙm#6ҡWd��{n�K�H��CnCo`y�НP,L�b��u(�RD�IiO�������YSoBBY�o?m_�=faP����Tx��0T�i�`��K"׭ xA�#;df'��q�.�zK����y���A2	����!�B�F���/�v�l��(P�5�[ rƦ�G7����`M9�|v�k�L���!�pEq-������{NGÀj�O<��U�L�q����>�f������e�����QX���g��0�z1L��lcߝ�#xH�{9.�0�֘7t��F���"ң�m�9ў���#_��7n���\5ep�{�t�R�ժ�y��|�{�2� 4V���<��֫�	��v�����۩:��`9� h��2��b�s�gW(�OP8[�&}N#0}v�����eп]�ñ >�F�9����׀r(�UEE�e^[�h���k��X�{PW�Z���P�����@����k���|O�1]me	�XIK?�+M�m§U>M�*O�Ue�p�ƴl���|5_�����7��'��I��,����nla�$V7b2oٯX�	{ٵ�L1U��ZB��e-�7[�Mfq��v��^���AC!�*���v�0�L��-~C_��A�EѰ���Zi9Ś%��vv糲-���B~�ǔݏiI�YfOץ�ɫ4K�-sZ"LBC/�k��o�4{�ǈ����#o~}� |~
_��3l$�%3S���T`�q�B�d#4�@�����&�\A�vؙ����:�h�[�\�G��	�+9�B��R���%	��q�����j<%�������id��L#ɞ��	���eQ�گ��'�H���Þ��>vP�̢�xz@,]��| kg�
���@����E?X+�?�<7}�0��!�c�"�䰀�:����`zY��� �r��2ҷ yݴ���q�����O�L�)O\n�*��;8�gm�j�D�EBW>e^�hT��V�u�g�}A �c�u�J�%�=��GlZ�e"��F?� ��y��6rI�5
��y�
O����Qvʭ��{4���? �E"�6��~#H���v�gj�k�<�i8t� ,\�DxPd�ޕ�u�k!c��Wa�Z��4)��F��[^>D�9�bњ�Y0�5̔����1@*��g�5���:�1�;n�nĴ��װ�覱�,.^]�yN�B2p$"�݁L���gNߊL�A�� G��6�N���s�ۼ��d��W���S��}j'U)p��؅~��~Y��$�W!�_z�:/W�
^.�Q���t��Ǫ`��r ׸Db$4�k�����	�����`ݝ��M�	�&*�|�Db[�'��?<#��&�	č�-p��|ŁKU�����4��pw�T\�����]"�t�Z^��@{�(�Æ$�oi�C4�+O�۳*��.ٓ44�
�����3g����ڬ9(����|��`�ѫ���@�p�X[c(�F���,h�eh2 6W�h��8A@���I�J�ֳ���;^Ǖ�Mo�(��~�\;H�]ɁU�T8C�\�by/As�5���Wp}�s6���(���$��j�!$\p3��U��X	zY�o#D�h��`�=�m���M���T��-�@7�{\�}��5�?�ˌ�Y�Yh���\��1^U��=��*����Y'���k�]K�e���F����:����rN��Q�R����2�&���
�B\�C����.�����ut}6�Io�a-aj$�ӖX��{�����"�ÎW���6��Z�m�F~J��!m�T8G�/�!�eU+]'!�����I�Ωet�*�Kd�=�zK�GW���p}>T;MQ�S0n]q٧�E.�h��ٍɩ�)Y�r�MD�YA�u��
U���� 䄍�Ƶo��x�d����$Oct�ܺʞ�w��4:%A�KJ����\�MW���
�K���Q L��&(90T`l��@S�33'zE
��[���8���l�.U��mzE3��	�ׯ煴3��Hq��$3I^|����u�����g�"����IM
2̏�/�.�c�r"��:�UsUܟ���}4F��P������ޅK!z�W���\�6�F-\	���G��6*�Z���=�p����/-q�O!�2WĀf�7k���&{��0 �FEvL��l@�OGi�JL����ck�a�ݤ�`�¾����OH�`X�(����X?M��������H�έ*f�}jy�r����	����^tQf<�\��~�U�P�:� ��� ���PR�*%��}bc��m���ň!=
]�ےg��v$�����9CG/��՚��TFdM��fE�8G��H1��N�(^Q@z��i3'#��3���B-�c�F��bL�ҍ�^n��d ������j��?�\�t�Cc\C�l����h}q�´�s�b�7�_�ö�^�x(̅���V�_Fc�fr#��%��>'��%IL�n�Mt�Bⶀ�����}c�]�b{0�������I�yh�fW�׶��ְ�|䂠Tӗ���%�
m���[�>�i<-D�b�*�O�'VT2/�����K�������7����0��YT�71uά�Rgܕ�AE�x�J]]-����x9W�Gm@��	r�.揟w���G)����9�	T$��7��׼���\�5����x)�
]TGB�"ch����D�$�m���x%wb�d��{�SF4�p2�`9ǎ�;!|�E,�e\t���ЫT�Xֳ~�R��0v�S���gb���	�E�&	�j5�� �ф��/���ٕ��3IY���գ�Z��;����R���@���D�nH�~N]/���'ڴ��ǤrF�J�K
�!Ri��E�}z�C��s��D���۞�:��>��˔O-�W(��o�~$�y"A �W`���v]�t˫��Kd�8���}�X�j�<֌%X�k�:�4!=���A�<� ��Ը� 2��W<���ޕ�,8����Gk�Z"$\�2x_pݞgﱂ/Դ������nJ�Ӊ7��������Xh+ӳ5�0#>D��EGr�#=b7<���D�Ut��VװA�eB�qG�ܜ6�P-w��[��k�B���ծ`�>��8���IC���p���3�u'��Q\Pp ��$�������$�P�w^����$M�F�ap=��l�͠�#XH��) <����;�B�u9(P��\�)'+D��1 �:5Q�L�+v�bf��"����^7��8�v�+�Z�3���Tk�rYUF@� ��>�X��@��F�b��<Aה^��-=�&�s�k�[�n����/6�M��!#��h�0�@ػ�h�=b�a�9PYX��^��?�u�R�k��A��Ԍ���[^o������çp�J������{�`��2;�E�<�vе]O����7*�E�?�;�1��L&y_2=Ă,��%eD��c̱��)���5���r�\�rq3d�l�
��$C2�`������ ��Ĳ�x�W؈��=���u	x�KG��:�^m~�f���2���sZ�:��%4x��~�pL飹�����N��=}���c��η���#��O�����3��Fv��D!,>��p6L6dt����A�ߗ�	�R�D��xuJN�dg�<�2���O=9��zt��d��5�V� X'����55��	\:<M�`!�S�w�c(�TP�0�,j�����`�6.ǀCY}�-"�A�<TY�����N�����*C��<�g�z��S�k��;��䭿T� v֊%Ϯbڙ��Z��������T���bw� �20\��of@�EI��Ds���N ��!�@��+�T�fq�Ҹ�9Ӧq����Z��Ě�Md]�:}���Ia:?���� ��W��s l����N7>f�Z�9K�օ��������s�0��R�V
�0��&+ �.�U��~(�����-�R���PG���[x�9�+�֯@2V�T�����5;����d 5�c���C�7�t�{d�޵�F�Kۜۓt�٣� ����K���&��MG��J��qXw
n⎲���]r�*��vl�D��m|��${�r7BfQ5#FTmwL�+���}O��e��b�n7utb�Kkl�hY:c��=�nB{�����H�� 5P�S�������%�0���H�H�L\ǌ���I��S����DH�oµ��z1��1�B�9������w�'�H�~���&�����r�%-B�B�U���N�z6��_���D��1��9�G���S�k^g`�T�S��P����ʁ0���Vb�qv���<�\��/�~ހQ01ҡ��e:ny���kљ���>%?A���p
~+�g�$�$�{˚�J�&8�pG��|�����|�T􄟫�V��=0�2��:�W����f�(\�6��T����R�RxJ��ڰ!�Ni�7ج��J:O�#4�Awmw:=�K�:2]5?�]�O�>h��:��C�ҭ��-�V�/�{b��t�h@�=���@}��bׁ�%}�8댰�ڭ��ƒ�#E���Fm���s��/�3c��O�ڈ0O4��*1x��i����8�w�,�l�&�o�8�N;�
j�V9$>��?��P��O8i��dy�0Z��9�	c~<��y�M�$-�� C��X ��ܼ�i�(o�:���9M��4ƞ���R��I�@�G80��h�:��1��ȩ譋�8�sfe��ݠ�Ġ��;#��{5F� sɬ�B��s���Z�(zI�x�g��˯$�%��8�>_���b�>R�a���K��x� B�6T� �'��ZI��y[�	��[ R)Q�z��l��;�R��GBdio6��ވ�̔Z�%���n�Oy:��fO�	�1H��o���gi"�T�P���K�_B.;�>�i}n�h|)��߰���w#/w��<���D���^���Xˁ��z��a�>������4�ҀG	�A��2���<��Y�z�pr[t�ۻ� /줦#e�#?�8֬}�{l#hB��.
��3�o��X��h[�7�_�0]��J~ ԟ�D�/t�c��1��2 �V7;�yܳ�����Z��+}����k��Nf4����{��\�e*ڞ_p0�����T�!�^��Pн�+P��b� _���0g� ��ћ�Y�$��}ԌJ8�w���
|FkH���ˮMv�nبB��C��i�&ײ-��@�_ϫ3���\V��zCup�����L��'�@�a���)�p��E�Wދ.t,�Чc:h�v0h��Y�
�q/f���W��Ң��i�V���)sR~����y��޵�;x��_5�r�#<1�&����LO�j O�'��"����K���Q���itHT�[)���X�Һ8��}�R�{�@����O���Kh7?�~�߾f�82E[I�)�/1/�	4��B����%U�V����c#�&�Nv����Vg+2���_�Q�����m=قJ��n���(S��o?�0CD�n���}Z�d_��KЯ �}��?�m����o]�]ۙ/�=��w�������D�hV,��^1�O�	�D{��"����x��0�������('
3m�����Oٓ��ay%82[�s]nh6n����
�Lҧ% 񨴠�u�[(F�v�Puڢ)o��J�Ӄ��	#��T� �l_��鲟�qY�R�zo� ���z8��ps��K
�T٫Q5��pS������nH5�/|�ĳZW��}<�0�h�(ϩ����F�$����k��ʦEGKb�bd�����t�WMX'@��T�t u� &idB��+~pU����n�Y�v�_%MM���*9�s1LpY����\4�񇢂_[eg�g�2�p�[�gKr{z�Y��|��`cH���WF��mb>�8&'R����u�a�Pb
�=��% I�W<��w�)�3}�P�rߒJ�h�kGg�:���p�û�){J�6DG��_Ӥ��::  �!�/�� `3��Pǣ�C+�W��ݭa���Xq�����4��B%
[��Fo��ۺ�i��H؅�H-�TIKod��\8�2G��AP���)���D��PR1��b���@-1l������g%>��Y����Z�d�5��8�Ɣ5鐁��?ov[����'�ܶ��b�9����o�+�$�Y"��D�d�(it��Z���I����^��!||�z��\��>�Z�xTdP�9��)Q?m��L�뇻�I��E�r�;V��� ���L��y�$Ȩ�V.����Iۗ k�4-�7����8T� ��YV� o�%]�|�ͦ��r$V��
�8�fF�N�͋g)�w�;��/	�ܻ�t���[6��r}���9�]��~]W��3�CKU�!�߸�^ؼ��S��2TZ�IK#V1R�1�nv��-��[Je~�\=;����B?���	8�'��+QWK�/#~�!4��|mb�-�A�����p���ލ�<�GL�2�����sXS�t��*�Z[�l�?�W�~u��ⱻ��LWHvdW���`В��a��>qH#�R���x��8�IH�n��
�s����>y೓���PX)D[h�2�5=�A�/"K�(&�8O��c{�+�KX�Im�_��!!�)e_s0�έ��E�{��:�
(��qUcOTW?	���.��1��{(G��Ӕ��`��==�W���	C�].� L4��_3ׄ��]Rw�$���s�hWA�����B܂]��e)r�g�T��Q��OY��3��ָ�g���&D�XS� �3r��?ř=�����,db�r��"�U�q⓬�D-���d�Ĉ��n4dL�m����؇9I����A���i�sk�	V>�X*���J`P�Ʈ�>�_�,��#�S�\T�N.MJ���O=�N
�F�h�F�!�k�@��Rơ����/��ԇ-��}G&V\�p����,}��@�1����dZ��]ФA�k]�9���������Ev�/}6�1Q㒿�j�ҝKǃ�4�0�p>�RO�t�{ �����;���'�Z��ߗ\YyX�s�>ƒŭ6�_����x��%�C��,}�#,ax����g3�yA����@
�ܦ�h�ЌUmÉ��,X!�������>����s����rX�n#���g���"J�$\���X�#ZΠe�I�������i��4^� �5����������;����_z]�cTf�C�AR�h8s8%��dRzV�v��'A����l*�pq{%S��,�B-�Ǐ��&ڍ����"DX�e�χ�h��UOE*8��3l%��Қ����'�3��g�� <�/���+��H�|��n���Q���I�;��:Z�C�c俢�B����<&/�׎-s�Gl-��̥��W1z��&#�i{�nE�ea�r?��i~��;YM���	 Yi�xď3|O�G��r��4#��_(l��*�ڙ����ʃ�3}��xO J�H"�ܴa�1�s]�3R2@�_�`v�=�C��a�ӏ�첰N�9���U,f��;�9$q�L�h�� �z���T^�������ԅ"��kzLsR�����}��A���ӵ�7���DKy�[�I7J��Fh�"	b�w�0(pmQܩ�\ԸK������`k�Iց�f�ZeV"��ӫ�<�r����2u�����vKo/.���\�1H״ܵ�)-ʢ�����p`��Ud�7���mGe�����-�H�8��G!.@�XK`7y?IfS�v$�3�쓞���Jk���z+N�����}u�KJ��ļ#�n�V�{ɠ���3������u��	��@?tL[^Bl�t�qs���Z�JX��d�针& ��6�K�K�	4x�r?���E5_TI�lJ������?=uN5ئ�U|��jvp���aS=�H�Ic"V�J��g�m��Y?�X�YeO�	Ž����5�<��U�~�.�2� }B�d�A�!��)*��zC�t������JqS��)�n/� ��]��:�o�1� x~�*������{�K� �
�c�+�!:���'�\��2��]�̉�����K�(i?�@��xi�A$��$��*{��|�@~�,��ĥ��S3�(�\C��b|�d��Oc��5�
�f�	��2y���VP��,$�� N+���@z���_%���-�OlW�:��2/�e�,�L��?�g���p�.O��7=��-�a�/Y}���帆\���~d=U�[�s��h�'L�)+�y3�������@I��`W�P;λY$cv�^u! �E;��e����Ý���7�5�m�y{*����ir��Z���8�1�*�ص?]�"����T+��*i��b��6�����D�~�������ѭC~2n4�
�
כW V�p�wʅ <��L�%��k��-��hrKe���¦8�����v�=6z��w}��<r�?���pc��T# �Qp����:w�IL^�(㼡|_�
 ����z9��b��]8�G�p,��銊��e8ǭ��Iۂv��`��k�PgDBz޻�
�b�o%�I�՜A���Q��ʣ��JSqx7��uC֯|֑~xO�r(��e˖V�Tܯ`��u۸��=q�f��X�@�c�X�}���O�P�5R��M��t	/PgSiV��6�=�4~P�F�h��q�Y��w��x�c��Q9��=[N�p��,zӞc�/��M�ٞ7�K��S�ڭH<S���_��klzX����������=6�ibg�=���lbdLk5O@�(yI�9�9#��9_t������R�W{2�q,�S�w�(����T���К�Ϣ�5w�F����W���x�M%Ս���_�s���2�p�|ٻ�WE��;:�ep��z"�.�)��,��ʆ2S�D���H�V3�ُ'�q,-	�����/jإ��6ץx6-ty�8b�7SXA�#m����7Y�B�/<)�pv]$�_7��8_�D׉�,�Z�)H�S�ـ���}�[P������t� �K�X=640����kٔ	������RC��ME*u������X�b�8i"G��eq�SCJ#���|x�0Uv'�F\��KA�mm���zm!�o@��f�
�I9}��Ķ�y�35p���T��Ȟ1�qbc��sI���p,�'B*�Rq$>ٴM@�Y6�l��j0�%cN���$ex�1H��(<AH��Ƃlנ�
��� ��:���ĖrUi����+����5���K=OF���1�q�7zSc�C�TCi K��Lͨ�f;�f���A/|�;ߙ'���KSe������,��P�K�$u�����"�����z�(�[,f�M%�qD��=@��©���γ�L=��*��;�Z�"4��ru��\pL���W��q�����%�������sR�Tm�t��nB�ue3ᓁ/�"V�=��������o����Ьu})@�_��f��ve$������r�|{me�b:%+�k*��.ߍm���Y"�ţ��x�k������%\yYS�|;
	�&��\��ʖ'+9�N	�vf��L�F�\��X
���fj��Aµ4��%i�������ܙ�4KS����,�y�aC%��2F�.�HYj�{v�w��c݌���f��xQ�G�'J�~W�ӟGe�Ǝ���f�}�NƸ�z�ߣ6o�ɲ�x�b6:U��}��l�%k���2���wP�'G{�<���6�X���ŜMv������>C������5F]��D&�UԌ;�9��;Q~�u�P�A�s�+5@W�r���b�_EEFڀ=�Qr�S]����S�T��E�"o�[*���t
�Q$�^=��\�Kܭ�Y^�� ��LD���@��V�B�����q���i��j ��$��T���Ч(ؼ�w��n0�&d�H��:�Q���I¾|aO�NrP�U�ܦT̪�~GE������n���$�x~�W+�r���0���㈱Wl
�\��FA
�p���J�RKe���c��f�v�+�P1����|�Q�!�#�Qx8�R�sܗH#�'��������k7��Y��5��mx��T�#�����Y�͋�7{���~�q�4�� �75><��<�I����E|�=��v���o{�N�q�8���|�ݹ��Yv�RXN��+$�ܙAF� <���"�lb�JȄ�� =d�b�_;p5~���ҝZ{�E����	)=A����ڵ��G��Q��}�3!䁫� �7�d�������ߙ>2��:���v�l��G���y�ɾ��/���W93�*2�E�D�W3=.�H3�eg�p���W�[Rmi���+�|�G��@�@���ky�pF�
�V@a-/�}|-Ht�k�C�Op����Ʃ�I/�'�� I�d�MW-ʘ)�����*�.S���q<��)�r�t*�������'�x�ߺ^K��YLє}A������X��ҭNeַ=�~���wJ:ӄgn�^����Rx���sx74Z�v*�K�Z�
ԯv�Xq�w�q��k��:�1c�g ����؟ ����L2�2�Oϙ��d$�±]�4����|<L"�?i��>�nߋQ�Fo�A�L��j���=�F<�CH Y�1�}��*��lNyH�=*X\kv�Q�A$��rH+�0�x��^�2fE�dN���{0o��v�Y�!y;������IDC#Gsl�y&����Rmy�r��iC�Q-�-����ۉ4ZS�>ǰ~�*!�&! ��H���Y���(����H�����Ł��J'7�?d;8@�w�dµ�/̙$$W�`�}kH�?U���FS�0���oMj��蕘9@Cβ&�����E�3��ŝ�`�+�QB�¬����I&9R<;�����^�6��g�q-���+������
< =�55��&��-6j1�s�ɋ��v`4�9M�
�O1�!��~�i�F�q	�Tש�Fu��J'ϒc�m�����i�5�ԪX�~n%̜�no��W�&6<�u�饜����L�R���v=j W��7��fG�XE �҅DR��<��`e1ܙJGY-�Aؑ�'�%�����{ +c�]xbu1 ��+j(��΢�	��X��qj�e>�E-��Jx�� �b��y���O��[�էAAA�[�y��v����rh����A{~]���/�? c�W� 볠�8�g�\�ڽ�c8z�\5�69 YԌT�\~�:;ˋ6�2�SZS�i!�3�D�@�S��aJ.���Aя��R����V
�|��p�Ҍxy���	��?aX��Iy��u}j�I��o�M�a.ӛ>��oN���6J@m�s���5R��x��m��&p�O�j�c��?{�'�� 
��"��Ho&��O8�7��a��G�k
6��;�{9�kɉ�
�ʴ0bb�i?-�ۗn�:�N�|7�[X�LҘ@�\K������ӑ�B�b���g��t��6��^��@��:U����N�8b��c�3/
� ��9^����$T~O ��(�ă��Ik[e�>'��ۗ%�Tx���g����&����iv(W$��ا����t�k=�P�@'-�>�QX6#�t�ժ	c�2�u����|ﾡ������y�s@B��)�RR8�����%C���Tc��zE�T��}�}��L'��{0�����(�lE>��_��a1��u�S��1��{6��,X?zϵy��YO�R�P{��G|��{A����S�	d4{��_�H��\	�OE���K�'�s*^ֵ�gޟ<@���W��<�"��ґ�%(�Ȭ��v��+�t\��F�;�{Ϡ!�;,�=E
r�Ṯ��z�!��Kl�)�=Q��쪅c��^3��_�� �JS-���l��ֱ��*��ӡ^��i|3{ �z;�����:��&�d�xY��b �O��tRS��,�φd*0�����;a�sib��[�hG��1C�: 7�A����W8X^�ҵܭ@8�U�14qd��+�d�6���5/����.�b��߷_�1}��6�Y��7�Sý�Zצd���·/ڼ�e?�>��	�f�x鯉�@3Ye��0N��FE8�(�r��>Z�`��g[.�ģ�����b�T�FR@�=�S(w_y���C�YtM��$Crx�E$�!,'�^�\���%�o�݈��s2 bv�z"�����y��(���爾�'ͯ�T1����&�5�� �;�߻���Nʃ���Xa��g[���Ep��sT��-�u�&64��u�(dm��4�'��!A*B)���R�;l�`B:i�[�־���K���fy1'�P��{�i��1�)�ύ{m�`i�r�2#��}���5\�Y�����ǜ�2/�4���n�R�|�"��ۗ�U�yجЉ��pX�5DPx8�H1'a���<�>a'Eс8O=�{�u�:�Z���L��e��[`��N�V���H�+8ݿ.�6��h�����N�P�6�K�O���ٶşu��V��ᔎ�w����j���7�ЅݱeU�}P-ɨ��]3a���qݎ�1 �*��n�I�P��"���%Ծ���e_�o�����x�ъ���������1�D�?��<(<�L��8�� F�Q������&�PF��O���-���ڤ�8&�h��'X��.�:Pݬz2�{�w��x�.���32>sZ��u//�y�	��D�p�ς�����q��ζ�}dV1�mC& J�a�����2[ � ]�Z|{Nl^2`%�+�7ߎze��V�(��� (����}DV9ƚ_���ʂ�_葶:^�:!���!�.�W��;���Ը�x�X�를�_�S2�	�u������A��.�� ��$<����,�*ń��>�hNg�~"8ryG��-F���9�ĜI��t���	�u�aGo'Ly��7�&,��(퓫�3�i�T1��Ȓ�?<i�U!��"�G3���F����y��ڦP~���i=��2��W}P�.��e�4V����&U�@9f�^u�H>9����||�ek5�vF�w���)O^�u�,�W]R8�����*��������k�$�O�����1���oL���?�~C�墌=�h�GW�ܸ7%^�,�Ijx��P����}d���E���r��I@s�N�f��o'�ۥXN�	0��~#|�:6��k�E5�����d�9�X�o���v�}���s0��a:UUO�O�1��ڳ�l�N��3�`�7
Q�9/=G&�Rql�zx��e�g�q�乧#�94���j�Rg��VIQ`���s��W�*xZ@8؍=F�x��HՖ6�r
6���s�s���2wF͇�+�\��m�'2�;O
D��:�=ŕсx��N�|y]��2;�o
�J��#������9\L��[8�EG��$�D�����'v[�y�&ڱ�a/��.��CA	y���s���Zk!�c���ѻ'˜&��~�6�@4����T��罵��#�u �<;R��?��Q���,�_�}1iE�/��i��뎹Ƀ��E�º�U#7�S9��~7�mO�
g��@��3M��Yj	a�^�C!YKm����w�\��q�Y�y���T����iKN�d�n�����Pٚ���O���Ze[���yr�-�m��S8���s0���W�|��6��h�*�׷�F ��s�� ��G��ۆ���)�~Mw$	ov=�o�F��TW	:�D���u���sޤ� �M� 8�^���> �$�?'���mܛQTA�X����-fwi`���[� %�FdԨ�0��*�څ� ]�1U�t߫Z��ۂ��p�\)E ���j�R��HU�����*iG5$������)��_m��C�]C�rO��J�d���N} �޴����^*,���<sU��pv��J8�O3��u�m���9����(A��f$8ܿ�
�����NM���=|�&���8�$c��XX�|���X��A�m�)�)�J�&�[�-�f�}"��	>l��,��B�1�
���؎�]����W�*_���N�W◭]�`�I���u�P٪��Ҟ��\�a�vx��S��<6[��u�B���;���u�j�U�{�� �X-'A��b�|�|]����ɢx�h���G�~,3�ϑ����t��#�f
�qm(��2�B帥q�3kͥCϏ�GK�}����=�q?�5+��?��~e*E%NS8 7��A1����qds1�7�����}��J(8�e1�zl�gn�������t�K�f���4�*|y���.HP��՛t�ɓ�D ��T1нrɡ�W����3珯;汀m �����(�S1i�X	g�������1rX���+I@���4�.�{��{�c�!"좋e��껈����G�f�y�&�Nh��)`K� �d5jh��3���=�h\��C/������Gu��W�`�!�L�ᨲ�?}��R.%DM�>�9�E��o�1�b�����{K�B���0�F�7�!��N�N�u�"��ؚ���y	?*�A�(�3�1�ގ$�-��o��嫴5!=��mIݾ\�.��blWȁc�:L�R��*uZ�Pe�w���fϥ�����.{���B��kjtr�S_�g�yk� �X76S���|gT䰻'-U�
j��0�{��F��x�?�`>>�͑L�\��m�. �Ż�%^��W�	��p�+r��-1ŲY-���7��K�PI�*Gj��e�؄�l=R��v s����e�i����5J
B���b�t����F+迬�z�E��fg��%K�ФK���t
�c6�/+Ad�#!G�[�ǵ#
j��mo��,�P��#Ā\���$\�IT��k8�i	8�U �n�4BP�-(m
�2c�{Px�)5ai}o3?Pb(M`&����{�s�1�:%���iB�P��1�(l�N�i Tz=0؜�A
/��Z�^�%w�*!ʝ�9�<�M�E,ă?ҝ3F�Gpc\��z�6��!b�� $�Z�t~q�>����M��ί��n����K����ʨP�
.�p!�L6���Fs�8в�>���{�6�@�
�n��g5+�w ��ȓ4I����Q��	�}�*p�&�EZ��t�������W�֋o�ʯ�F�UoLa`�#53c_(#W���Ʈ�����qW��G�D�M���S|��eb��m|Ft�q-P�JU�91�*�'�+)���-N�=��|�c�z�}2�l��Mm}U�w� 	6��9R�.k���:�W �6j��GE���u�LA���i͘ϋ��v�w�Fs��k�専H�����^���d�:S*�8CGo۵���Տ�n�뇚��9�l�N�S+Oq^�I��a��z>���>�X��Yb��W�š��8#kz�����`my?�S�+������gÌ�ea���"�8U�ZV�a>��{&��](��M�RŪ�[
�|N�M�K:�y�hq(v��f#!.��/B@!��Yx���]ZEXee_���W�a��ᕎ�/;t���>�aO���3�Ee�ծ#����W�u7U¹,���U6�K��yo|�,ԼN�
%�[��5S��9 2��czt��)�{�33��8U���W|��m��4�a՜-N�k�����l�Ex�����>���1�p�㸂fRX�'-��0u�x�	QHp�e�;��
(�d�'H6�p½DK�U��MC�&�)E]Y�NB�4c=�=7�=�ڸ�"Ţ����h�cLG��d�b ��.�1���^���<����n)��`k�2�	Hf�
��5�BC[��b���dX=��G� �����Ϡ�m#�^
4Mk��%�T����e?ݎft�8}��$�O��n��"���	S!*�	��;|C�-���EƸٳ����=��ݿ��N��s�1����#�Q�b$k�6k1�{S���B9t�L������"�y�ˡ�0q�1ȹxh�AH�����m r����X����T㹯�_3Hn��8l%$f;xj���<��RS�RT^��F)��a�g��]�����VG��`��7�>&��b�g����:n�}TX�B[T~l���
mXdk<%�o�D��E	���)��ux��_U6&�rao�N��̤^��6z��+�4a�I ��Z��U~�q�@����+5Y�������W�xpE<v G�ꋘ��i�g�1�*�����z�`���t��t�	� \:���S�򐺀����a��!��b�����G�HVܦ�)��1H1�~fd�����z�w&x�Ӑ���j��7*��;�^箋�%��&�WɄD!��Y獭�A�.:�)&��^����qx�?�eߎR-΋�ֺ���_5�i���DNO7�B�Gxb�hiF��gG�hWb���`����'`��m.��Z��ZF0�v����n\�Z�P����رv�JCU)�A�����X!h��?�^�*`�jkU�e�v�m�+y�΅��E>ǚa=�3F<�G����tɱ�#&���9�G?��&x%��<~�q��	�u���W�/��w �{/\�n��diC�[\,E��z��-&m!JI&�xmm�Ԕ��s���&�gf#���')� ~�:���c|��7��G�Ž�e�t��H$�#ݕ�ж����Y|^[�}���̣�M'�� n�q���U��j�VF�GM�,� ��]&噬{^N@�� �u滛�X�$�����+A��I���cL����
�`�o�{Ax�����F�ܒ��@��5?9��-:X�,85y�Q�JЗ��ݾ��K)����X�1��s�����;Y�YH�������&�D�3�v�V��c�G�bJx�?��K.��e�d�Y���+z����v����a����4�0��}H��[$]��]���_�|�M��Ʉ���%q�K4�Y�n+��Z��t��o����fAK�0���red�q��=@`�s�_�+���<o��K �FAhF�Z8�i��/�'E,;��2O.#":7��<��X����Б��vwE��X�H��tXb����
#�EUZ��F�x��jk�6���
̮�U�1u�W.��5c��2�4��)��7�"�a���U�i
G����(�7jĥ�M�����������{f�"dȐ��4�
vL��,>a�Y� Ht�[y���y�c���q����f&"g�rB�`��� �S5�.�|������A &$@�Ώ�XG�(�4O�L�l���f��q`�U�_{\�����fm�NCDlr���~�!��@(��#UN�4��JFE�|��uR�y��%�s3��>���-~{�A��Z��H��/t� ��oQ���I?zCM��Ĉ�5�T0��oc<��˸�s��+W׽OO���D�����b^�'Zӣ���j�7IV�bH��J���$b䍐ɣ�De��l�5'��_9a�~J�e�Ogq�2�Mu��A+�Ҭ�X��N+/'/C��>��ե�=L֓��:xklr�'[���*���\���������Y�3�n�l��[g/i�Y.�F�J
^�ה�4/丬�J(��l�9��)�k�0^��A6���es@$>$�5��UZ�=(��5�,r-MG�����a��,M��s��s�`�������7N�]���ר��e����'F��Y�X��.<_��՚�w��I#�b[<�C��	�0/<2Ԛ8>�1�_�̭v�*|�G�d1�إ�N-|E��q+�կi`7�\{MSG���!�V���:d�1 �\vFy&Idr�#t�V�#"�)E�;M��u�{ե����z+K��WIW�,T���(���r���5�_�<֫OԔ}��\�0�>�W�����)9�fq�$B�)[�}�������R�����e��� 3GIO��c\�!Қ����T��ޜ���2If�6x���⌠(C!���G�!_<��XVb^
�f�[�@ye�cE�y�oQ�(�D��1�y�����y埕�o{��"�$�(tt`+�0'��