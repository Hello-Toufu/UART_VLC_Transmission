��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��P��=:� ����(�)3�� 5����l]0�ك[�Y�qޡ�(���fZ��#b�}a�3�
>cO��o�LW��4�C���(C��&{��"�v11#/I�&�)�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_��r��)����%|j��)����kMd{'��_�$�iC���ff܀���o��|��y�Zt7�ׄ�'抰�i�o"���MQi�n$�w�3,�
�r�%l P��l|�M�0a�ha��n������|��!<q�Ф���QG�M���ȝh��t�)�����������=�J>��(�� ̳ݏ�����&Q��X��4��(�PC�F��\�!pP��tO���"�q��������81U�8����=�A�\�9�Ȅ�'�if�ŦizvTf�������R�]n��u�?�r��y^FO�����5%��B�ݹ��>V�8�����5=�{��;P꤃��A6m�W�%�ڷG���~]���n'ʢ7&\�c�>�@V(nԯ�.���~����ʏ�E%���(�Ǥ8�g֩<ȁ���M/(�`X�&)�X�
Q������f d��2>Rt���n�W��1[]�(X��a�e�,��B.Vd��e)��Lk��A���^��y�	�Ѧ���(a�tYhѸ�~gF�g�����$5=7,ʾQ n�/Y@��1q��ȡ�K��΋VSPU{�P78�R�0 �Z��C &�Ժ�h �=[KL��E/�4���LC��$��H��)����Z�p�/����mƒ���H-�q������v�����|��05m�E=k��AD��ړԍ}��