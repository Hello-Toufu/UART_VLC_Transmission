��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_��Ջ
i�xH�	��P����U4��  ���v����P,�u��{��?w�B�U�0���;G�v?��l��Z4�"M�Κ�Sq;F��(lk�]V'Ӭ�'���r@k�H�86K}�Z��Ç%pw�`4�:/Ζ}E����"��\-�nDܶZMv�J�O;H"�&<@y���p�1V�hR��¯@}��໦�M��f� h���^����zo�!�6�mX�7Ame�#�V�C�3���C[b=��.��rJK�Vtp�����)�κ�n��7ϴ��]�*�ⱜm�c����%���q�"��1�EA�������)ϐ��O1��z��4Ѳ�m�e+�U��O���V<oX����h�ާ.Q�0�}�� �=�(ȼ8Lx���U,�Q�^�ue�����9��<ۉ`k�0^>\mT*���9B��2z"�;]x�2v$��c<ȹ�i�簟��)L����C�fX���)v�L3(=E���R,Κ��fe+���o�ou��^��.tS��v7d�d���npp̈���y�.c dΏK���fC�ȘȗWu<�0��^��\9 ��bm&�������-�Յ�Ì�@�.q���,Y�Ǜ˕6��1=�������sE�Yz4_��j�!�q/']�É(�����&;M| ���	�j$�Nz%��`C��A�x%�3} �CJ7w��w�t�smw�.�F��Ӭ��� ������)/,����Dv�Qs���Sb\xF�!���	��M��Y�j߭VEF�=��,n��XF?~ή��ȅ�c
�hs*VL��7W�B�l>�W2M��M�6"���JI�>4��h��f����@���~a4��Ot'۴�,.A�}��L��,��牪�]��!����J2 �8C~����&�8B*(�9�8jQ�`'�-XB���$��^ߊ0R�8>,�ߧ�"ԅ��-5z��Y�U��VHg�z9b��䃰�;-�6�;��s�����}��D����X���S��5N�<��8_m`�֮K�@�~����̋�(ſ�$�O����Z���o���g>(E{�������O+�[�����tA��%d�mdԫ�+u�xЩ�wg�NbH�
�5��Dv��w�)&�M�G��=�Qï�H࿈�J^���D||�6���h��<R�|����cTA��~�\�>�-�:���	< �I#zWLQ�4�=�	�s��Qd?s�i(tޙx��Xf������Pz3���w���-xxS���əQz��qu�aFN)�8���C���d|�����yb~�j�@cz�s��EaTҕ��=�
�})=����Ϩ�F�߻x�q�
���V�%H���Z�|��y�4�e�.B�ל�i�&o��S���S^�F�h�~���H�'���%���6?�8�OmoP���.�����隀C�P�J�86�#_V�����]\pH��Ҷ'qyM�5��U�VY�t�������A?����r�B@�hB,�4��qSi�����#���eu���&�le0B�w��[�2Ic"a<)� �����/sk�m,�O�!��~#n�z�'s��K�8��UW�u u�g�BK-�]=�e>٘)����D�.�r�I�$��֦�Fx���"<a��yP���>P� �4<����C�J�2i�w_)+�/�HZ�#�CA�~��gO���X�
�+�LaKK�7.u�r�c�|���	
��4-R";(vò����HZ$�B(ݖ[��
�,`t�2gkp�e���>a�/����哊M*��Ws�.�j�� ^�[B G�y��^��]����/���.���Vj�sakʔ�t��F���X`:O($��="7����&Hf7���O�E�D�)���3�����Am��itGt-(��Q3�l��g�{J"���s�>Ft+}�|��}��E ~��}qI��Q�#N����|��C���I���D�q�-��w���}�x4|9&V�
�|�@�ҁ~0�,m�*$ ����1���Y��5���W��Q�H�}��sCN�%o�{��z��I��1D��@!�Tg=����Nn{��{)X�U��6�3Ma�X`�<JqG~�>��g� ��-\�?��s`�G�#���N�^n����a�i�	��Ӣ�B�,�_�°
��3v^v�2Q�h~��-ݍP�ц�:�a֬�;ڴ�R��Pk��iH�H��c�هr*�<�|՘����HN.b��������n����C��n����2�kԄq�Ԍ�Y �'�y(����G:��Cp@�*�5�ыŀ �!ԷJ�K�X�irHR6�kī�"W�N��3O?�=L�b�e��&o������6��ע|	ޢ�GկN�K�v|��1 gs�3��E�p��2�۲[_���͑��D��GG2؆��X:��
��i�>��طZW*cֺv�z�	���<������vIӂ�NJ�}���=$���x
��g��R�ҺEE{���[e��yI V�k��a��
'.G�_�6L$�]�DK��[P�}���e	0J<f�T3�9��Y�*��4F�Ǹ^u �D>k�-C�N�}E!��N1�G�G�6��bdm�E��ʏ���X*���S��]�t4���c�m��B�^Y�|T���ރ_���u��a�<�����y�o)��5J[h|����nB�c����ߦ2&a�6Ĭ���n�9�~����+��e�t/�/�z��L�;���b��dN���%N�5���W�b���mP"钼C�G}�c����f|����bQS����{��R�[Y����7OL��L�):|�<�\q�@CHǈ?��L؅��y�����pn��A^�e�w�{�]�ln��WÂB:�-� ܗk�W�˒�b�)��Y�]W�k'vK\w���kQ죭�0��j +�ҡ������/;匓����XTI��H�`����b�2ڬ�X��q�O6�s]J\��g	*ZL."fo�Y�U�܇K�t�䑾_$OŸ��32���T�B h7�*J��C����hFsZ a��c|��\I�K��\�Z͏T��A=��t����/�BH�F�����u%Ԫ
��ӬR�G�9촇|k�w��U�Q�R��PaӰE΢�N\�w��W���G����i�����oɔ8�qP��F�_�p��wH��g��k�W�	N/D"����&\(l�ӁƢcL����_\Iڸc�S^Gǆ@�MO!V5��''\��K�*9��$7\ZKTՙ�򏉰�E�I� ��.��8�$D�����}=��[�LIVu�ô�p�
�w�������L�r���{����i+H��}}n���ҟ���𓪚&J�_ξ{l�p��$ fվ�É�F�&�X���vN����5���flr�@/����6e��i�L3ł���uW��H��ɞ)��y��Zމ�Kz:���s����2~T��E�GI�H�iS��6�~�%��;z�����P��ï�j*��7�֠��TŴ�x�u��� ��z����Ro�;.F�%�\o�w~#C�w�qj'�DÙ�\�8Txر�/��r������8`@���Y�8������,$X�dD�o��v�d�J��]Wz�1�]�ꓤC`���<[ŉ�|ힻ^#��9Q[�|�k�<�LL�wd�ߟ��[�<P��ٰ�6��	���f��F���آ#O�ʭ�bd��=����ZJ�^1�Ӣ5�#���1U��_�������<�*�jp7MEG��Ua�%��ʜ��z�zL6��������ߤ�h<�٠��RB�.�9Pf	��M¯[��+¶�A6�[��?��T�l�)j(0�V����פ�q�ĸx�K���M�)͸�`���a���I�B�3�Ǽ?�x�0�mM+�Wf�nq@��.�` sJ��6�#3��t�k�i=%RLјܨO>��=�:F�=?�Si�8<f��Uf�kt���T	��,��5��@�h"��G��Fvr:ɇ"H�w#j+��w�,[Bba�[�-HMɢ�RD�S�?���H���\��\u�h�1��#Q��z:�жv��̣�;Ҁ� ט"1�}��8x�������N����D��?
�nPj��DO�t��t|HE��8��n�|��k �#k��yH/�����y�T���36U^�lR�B��~�w+߭tY�ë
�g��Q-�О2��=a�\04�'V�]�{n3�����:���C��@����û�2w�%��p�mҘu���\�r��E�)�bz�^�y-���\��x �b�Ó�O��}�3��
�%�����Sm���6F�ك�;����\1�k9�֨R��S������ł�
��Q��j@p9a��M��*�!��Sc�K+�C�8��>�{^gf�7��*�˥�� ���j��������UX���y��@��I�������,��:��ԡ��}�G�֠-)��'���0��8a~	؊a-`A�����	�mׁ̥�~HDH�~xI7�nJΔ�j�7 .c,�Vq��A��j�b��S\G�E��������Q��qf2K�|C��(�y��;�W1���,-�g1.�#Hd�N�4���X�������[]�2uPܿg?ׇ�`ĕ��
�;A�V�hZ6%XK2��;�����/)gjQ��ᵟ�%'_#�H t�
{n�L�����r�6v Q�>�b)"\�u]2����(l^h�bpP�)#1h�[��7wa��7���Y0oJ�T����z�y���zѐP0WN��SqJ|,�В�(�y�_Bc*oI�]	���S�>8�R�]Ճ�N�Sspn�i�����x�ư�u6�	����I���y���z�d�$�=�:x����!T@t���6.���Ȩd�
�߆wϨ܅��$�� ���Ń�Yf=@�\����l�,�oWg^
y���-�c���ż��m��@�>S����a �%��؃m�h��Y�%f1�E�srfK]gy���E!��3݃�]X�76��XH�zq�@�{�����~�ή_�B�ګ{��	�.'��B��������5_Y�� ��]���Xxċ���S˰� ��c�mm�>�Úc
o��k {IN�=���SԨ(E�&D�5��r�h�WI����W���J2�]χv�B�:MMW^�N���X�y�-��{�V޸j�q�N������h����8Xe����.��8�[�G�"+�u�N�dL%_�m�s����8�d�!�P���|\�3K�u�X�0��|��'��&�`+p�~��\�\a��4 Di�����!�ⒼH�N�3�ja�I�$�(�Y6�K���w2�r�He�}�r���\�p̕go�K���������ۮ�LH4ˬw�7�N"Si�^�s_{�1��]S<��-E�wv���4dIk�pC����Cm�"���MbI�*
� 5g����Wӈ{���+��E���ߒ��Z
ʁ�0�'�$A�����R�V�����〺@N������s\_rz���h6.�91�<���iYP	9����K8�D����8�������� �6����Q���),��Ҧ�N9����پ��=�_��+�@��D@`��^�[S���Am�����b���>'��
��	 �5�s�qS�
pHY_a����Z��of"�8���a`(#�l��	�er{��U|q�t���K���(��6 `�n�����,2H�-�3W�i��Ս �_���a7K��~}���r�m7z&�Df@)�Ŀ����^�p�Y�����!�"�������=���<] :�ޝQI�v���2��<:1����4���kUԻG����>�s��|�H�W��7�F�&��â���~XQ>��7�����p-�mĆ�0�B��tԉ4�;c���4�]z)�1�`�r�J���&m@멹ש+ �ug:�OAAb��w3��
�z>�ی�f��_-c��:eG88�o~��0Av=!NDZI
ܵ�R��tBf��f bTy�z��l�թ�-[��̡-�u�BUE&�BR�
�9��fKǒ�3z~�
����v�LH��]}�#� -Y�t��~Ȃg��k��cD�^5{Լ��P���9W�l����o���=Fчʱcֵ�1����� �م���� ��J.�˷P,j�ݳv%v��{M�����ɼ)���v�+G�d�
e��j�RLN�*���|��\mJ� ��x%U!!��.�ךr\&*	.0e��;�t�:�"j}mr���}�T�����9�W�A������y�]�4~w��u�R4�I8���U������
<�hQY���R�j��?y����qK��q$v2�KQrb�a�;O�V|e�$=����E@��`NC(^QD/is�U�rI �G�,o��P-0�g�D�����-����F�}�����kf��7��P�n�eV�3K�6M�$		�pN���%�(G�V}��XL�����gD~D�fV�a�J��:����,�\J�l�S ��,�޶J:����-e�)�	MJ��ܺ��24{��G��F����K pt���H0��]�v\�hҩ[��r�ݺCZ�&o�d�؎�E�߾���.崯�y��(N^R�g*FB8Y!/M��8G˻V_( V�+�88���=u)$Y(AMd �i��=؊>W9��5�~J�/Ub��ذi�l=���( �C��M�2���N�a!I��a<�8:_�S6��8LSc��I{�+O-�Z��k�����-2���Y�����P�}�BZ>��Y�KD]��2Du�@3oO"F��>ѥD$ek���ȁ�q@�V])y�+�fP��Q�b��]5���U�,�	 ��Q�F��$�K��Q<N�� җV8Wk؍Ab[%�B%+-Dз^sMy�T� wl�N�X��cH8��s��8#n��SA�4��{c����^y�-N��&��=@�M��[��X���hZ|����z��	"�mB�jw����~�A!�v�b���+�1�� ���f����EfR���ms��|��z �r��:�����=ԝ^�L.�P��DF]f,�3�8{)�5��r�yP�@�Ƭi=��0g��O"�Q��	��P{;�V�=T:\���,��6Zn4e�&�X�1�hn�$�r�-��;BE�V��%>oS�CL.��5�w�ٍ�����S�s$d!��,X�����O��E��] ���l�۠t�-�(�~զ������^[.�H4j��(�@ǽ�B�ZߓL������{�b�����Ֆ��O���.!��rv=�R#a�	:5�[_k$,`�|]c?�^0oLR�؈�!��1"���"�Q]�ށ~(��X.^*�Q�,d�ƤA�[�מ]ח��tDd�3h�hpH�~���W��g)ț���̡iv� �g�~ڿ����a"E�*p��I�Ԑ�_��g����ĦM�.�+m���ټ	x��W��?���x�1Ђr��ri:<�>F@�D���h^&����O5}3�9��a��w�ULLn����h��d�Oc�tݺ�y�f��H;#���gz�Kl����J)�)�M{�^ NiLs�x�����}Ez��\ۭ]�tm*o���-�M�H�e(=��	DI�����=CLꈂ���8}�<�?�wО��i3ǥ�;���虹{� �2%R%�Ҍ�q2ʪ�CR훵�o:����u�'\���E`��,F��Öi/�"¹��w��SM��5++���_�\tm=��\U����yː��;�`Bv]���W���8���)1����ӑ`�o#�u>nX��-��	0|�D?Ȓ��h�~�O��-{��n��A�%c:1����S(��x	�c.�G�����>~���+�����7�3v�.�o`�]W��e�� ��?�Bmc�	
.6�r௞�b#�!�eŔ�R+�N����TB��E�<B=@�h"�����vS�A�痮���d��FihvuK������;c���f-��ם���*РK��7�Db����c�;�!B�Ĺ�����T�53�s���v�5�t�Om��3;S�gl�^��f�KB�3$�ݑ
����ⓘ�T|����wL���d�s6��iL_z.=�u��&��}<W
-=RtxAhb��j�٦,7�V�6$A���e(ĔC:�� ����?�U��%|�<�V��6?�J���-#$J���_uN�����k�1;O�l[�jW�v�W8�wJ��?y5ߑv��?CY��VT���؊$�Z�>ᎆx�4��G�_۶83Z��t��/zE���,��PM�� �	��1J�7��0�Z�Ҵ�("ٛ�W��?("V���3�
a�\���_��;LZ��`nX��!�?� �E�M��'9���e��J3^*g�������|58Z7��A���}6 B�$|r	7�t�����k5Nm�hr������'~�q�/��q� �(ʎ��7�e�G��}\2`���̧������Q�H�W��纣Dq60l�Ǣw�
�/ل�ҭ᠏S��IK�������A�G�zZ�z���od�"C�0�ުI�ˬ�@ufN�+�NN���=����~=�KA�_�B�Dk�H�L�ܔ�<7�=S
��(�D����~�5�F}nToCCbF�~�m��'%CY��7tFN5Z_�`=�ry5�<�[�/�u(�ϞhM���=6`�
����4�kpюMl=�LB|���7�.�.E��;�trE;H�$�F��g;Eq������ڱ��L�ԝ���$��L6`�m��24dP�Ff,!0�H���m:.�Zw��"���f�o"����>�R%�Y��C��x�^	g0�����5rtĉ3��vv�5�g�4�3S9��m=Z�_�o�7H#tj9x#�i5g���ؗ9a�M�7k��F�C
,��J�Xֵ�2�̦��v�xa�f���L�I��~W�!
� ���(����25��9'e�a���B	�b��aa�T
�)"��ݽ�X�v�����K�^�������	��ԋ��%�#�%�����z҈��J��~9������	�6��w2��k�ۃק�&F@tOݨG�ٵm��4��I�&IK��X��S^��W/mjX���{{J�R$?Ȉ�3�s��؁ }�0�*�%FJԴ�z��æ/r������~�L�TA3�:ǎ���UL��?�$���]��W�z*s�}!�fG�������C���3��Q�k�U��*��V�ҡ����Pг3�n��^�8���L1r����t��?g���-	
pʆ�r�Ï�ˮ6pN'��i�Z�SrЂ��O'�����u��e�Ȑ��Rup%��VMʜ"���AVv�ST�+?�߃g�1������|�w�5���طI����U�]:İ�k���A�K�)\� 5�L�RR@}�v�+�Z�����xjU��itJzx���r��>K�Ŕ��
r+�M�YU��5_#HC�*�\��&��U?�͔�,��w�l���#��� )����������ʏ�/A�o�T�;G3護6�/�[x��!�ǮƙM��hk�ۗ���0���B�k<��p耪�?��=쀡��.�$�4$]���=���*8��˘9i��3MRD����|V��|듥�)f=��^H�#gӥc:ֆ�3���*6f-f�`� �$ߐ�dW��~a��&O��l:�:��Ypv��t�dzKpBY�홃C4�
���'��,c��D3oW�����yh�Wt�f!����i�^�SXM<8�L]ًt�`����F���{�d�]��ZM��Gkn�.�CQ���-����+V����0�`��fu�n��k���4��-��EB�0�rj��
�V�M��O{�2�p�N.��W�X�#��n+(\:��M��x���O�$<�F�3��$�kEm�ͩ�^n)Y��IO��$�ĿSl��(*���-���cbb����2�����Oj����i�h��<s�̕�Mв�vw+�*�n�Bo��JX����jYa����_E��z_̅̇58�I1��Ɲ�Td�)'2C^� ��ĿC�#f��/��.z�|x�&J~��D�L����Iv�}�]����<��P3�l���	�IԀ;1c���;�.�*N�����ѴQP|��a��k��=�I+��9��ω�սC�d����x�m���"��	��"������O���Q�R�@��o��ţ-L�}_�ni&�e�f��&ʞzN�Pm?<R��@�`�uڨ9A-���;��:�E#��VO�ug}��7r(pw��<��h/¡�\)�6���$ybNzt���d���@ev��>��S@����^��L.+'���|�T�#��:��"�W���:؊�pf��o��� 2��Ӕ�	�e�^M��`���@b@c���vwi&��Ս�i�2�4~8�/��$��v�w�-�L�#?[�GKA��M�ܰ(k>����ɻ��,,����KF�+�:�SV���=�=�*��ԣ5�?�5䒤n3�s��>���? ?���~��aޢK��,X���;��hG|��m�4��k�J���ŪkLvpl��0���$k߉?�����Fs�MqZ�8M�����Pw����!��L�y�n��D��m�f������' ����pmd������X#�׊lƇ_.uV�2�:��ͮ��r��4 �C�����F)A<郷\2�0ݛR_n(
}ÿmÎ�:�b�(bk�01&��kXb[p0zlCa���������%�ݱ� 9�M�A�)Q����G_@�n1N� x�%����Lc���>w;��{�p�����f�S=�4bi����������ʿ���a�Ǎ�]4Կ������c���/�^^k$��ā�QG�)�%Qq����ǚ�f�_��.�'�dBOKs��EK"N���	:���Q��WS�	n\��;Ii�\�q�k�G�ǥ�D��N��n���a-I�Tَ��̺scc�TI����1$�(���NGR��x�¹��{nYuvo2��=�B�L�\���B�MUX��5X�h^����k�j�@ώİa\�˖��So��/E�pk���fOe@�i���C��ɢe����l$ؒ�n߉h����-�����-"&�������q�#�S#�H�����u�����Z�x���nc8ֈjs�-�*�+��Z���m��z3}�D����m)����~��j��5x`8o���qb� �p싙��b�����I�A�U�IB8�c�=S=���Xĉ�>JF�l���Hy�l����r޲�A�C�Ӷm�Ǫ^��.	t��v$w�N7Ѹ��[��OQ�������/��u�+�=��I�J��P�
�WJLH�_ļ�����{��!��7p��%	�	V�Xn�B�YpE�&�#�s��-5�/��*��E�iy��Z��,�W�	N�<j838V�>���X����O����v�9.��eE{?��o'��$8$����#��(�*��Y��&�^��M|l�/0&�R .��ek[2+�VIZ&�U�'x�o�uM�ǲ�D��؈<�n�KVD9�u�ę�C!8Y�h�āo���=�y��C�HT6m���h�E0ڧ��E�9i���������pJ�K��~���W_�W����*�{dR߻��qWi�soo*0	�
�s��"��;E�49����V8�=�k���yv�p}���P������b`���%������mw���sb%tY{1^�W%�φ��97)��8���q�9�����Y�X�1�)&����J;���K>bʾ�N>E�YДю�ji�m��9�K��@gu���Y2ێt_}|����f�>�^-#�5^�C�P��g|���ɚ��8wH�}�]g6��s��uN�Gl{	M?$h��H�x �p[���u�3zҜ�~\��#�}�L˕����-<Ý�K> �,g���q�z���Di��{�ò��j�p7�k~��.iR�I50��rk�92M�
�D�RvRd��BG��Xc�h!{ʁ�V1�w�-�T�p޴��q��b������k6�	$���qɍ��2�7�\f��~a�U�`�qL"�@3K`[�h�&.����-o�E4`63�����ń�7����I���}�Ւ���l�	K�Z���y��Y�$v�x��j�Q�8��r_�Ѵ$���(Q�Ͼ�$@.��������YN�O�里�;Wd9��E��h: ��Q��Fb�jl�Ƈ>�FTڎx��D�>(%u�b��(b@��=�����J�=�_}�&}g� �|#������]>�T��b儁X�n��n�*{���e�x�1r�o�:<`Ou����5u�(Gf27.ы���Q�Ė���'���еad���:&�q�� �� �"[����9�"v�3��1���is�E��V�D���Vc�#5�ò&���ŮP�յW�6����T�e�7��<E/ĨK3����2�U��3zn@Kә��"8Mb ��H�Tx���S���_��p��D�W����{I���4|+�)�`�
�[��!J��T�#,F
���.Ş���|T��5˚Y!Wd��H����`-��.p;��G���7��$���P�&Ą�pk�� �Эw���r�l�Ֆ�
,3D܀�YP�`��Nş�5;	�XO��7#w>+�h�bUg�F��i��W��&����!C(-����+�U����pk���Q���4��$0�_AG)p$��8���L�ҭFd�M_=��@X�YH������,)�6��of:1���:PON�l�e|��ȱ!���ǀ��F៘�(��(�?7X��W�3�༬�y�b���@��#�y��r��B-�a<G>gIM�k3���J@:F�{ba5쯸S�S4km�b�eo|G×ҫ��`�4�����t)-7�sКxg�`���@�g'��oOJX������4Z
�,�@���K�ыPv���ېA�f�鑝]�Ћ�"�����0W��9��-�O�2Y�k+F�2G՗3 ��6 ǀ�F�P��gf�ईf��"�@�eL�7LbͬCO|���b3"�g��
;g� 'O�Z�Ր����e�i���R:P����:�#�@j]w�L,�"q2Կ�{�ֲ�(J&��0�@�CԒG�����۝SYe���I�T��E��l�iK�'�su��GB��w^y:WJz���$�uq������A0�h.?j��K�J ��tDd��Kw6�|�$^���ޭ��*O��}�\���p��3u8���7�����b.ɇ���|���6��n����-4e�ժ<hWL�����B������G4���&8��l_H|�n8��"�<*w̩��G�"��	�
�ʘ�&i�ۣ-��dW8�����TŔ>=�'F��!�!�or��D삧zaN(b��
�B�~�ͅ(��2�C1���~��!��3�����j�P�>��@:��AV-x�Y�1�Ox#X,�c�)��e�m<U�o0����|Q�@mh�^8��y��ˊ�?e�3�O����>ې\���XQ0����}�Ɵ,f��Όsh��v����c���m;�h�:t{Y�4}�[^^�7����I���v%n���Q�őN�^�i�#/&}l=�� ��	ܒ���J�̓A�aI)09ˁ,_���>�:X�b��z�d�B�_h�l�~ρ�T9��t°���D�𞠘������׋�Ϻ���yb>C�@���<�U~��f�0M
�B����R.�v��A!3H���⨟����-A�{_뫝 ��fn+z���'�IYY���b��W"R�������j�����q����;����}�HU||=�,���8��ug��V���P0�$6�Qܽ�>:��7�������g�f�\JF7������Ќ� �Pjk6�Sځ@)�R���-���sS�1�,�#��=�s7��G���u�!��:�1�و�\USX�ʹ���IU�A�IAL�_�YI�o�8E6��\&>�y4b%6���j��k�6�Х��Wv��
����G����[��������G�ƾ��F1:�b�~�]Vx���4\�Q���m��1���w�7j�t18��L@��>�z�~�1�p_%R��c��N�$ֽ��i۲�~'x�;�z�b�E�fOh����F��'�^��s���tx�%Q�=��H]��s�x�M(I�U��sdp��;
h����T6�����{��l�`����)U�w,�Z/O0"��0[���=�
ӱ�me�;a >T	��OG�?�w��~[�ДѶ_=|zO�4p�/<�#�����g����Tf�w�f��v�O:��t��k�"�G)��=@#�?�'KF2ϻ����GgnH=�¦j�Io1}8u����ls�RJ��6l�~.~~��� ��]���c��[�:�(�+
����P����*��t�9-���G�v���yb�q)���ܱ���z��cy�/��5U���b�/�6�_�FHc��N�番{_�������(���Ч�����韝��/b>h�=V,Ҧ�>�Ƿ�a�c���BI��	��h-�(b��C,�^� ��M!T���mPZ�_(�Aj ��oL�v�H��4�pK#���U8�\8���Ń��UF`&�"2?@Q���ݼ�91�}�2b�����E<��B/�#� ����v$�է�o�m�9�v,Ꝁ�:_RZ�O�h:�n ��Qx\�e6(��c�a1u(䵪��q�C���	wyS�����Δ>2�+$���I�]/"G�e�w��[�n�(+�~'0�ʔ�HHw@����B�y��P���c��Ƴ�-λ��)ӻ�/��a��w
�,��7xP����-d*�8�V>��4�`Bh�Q�G��4Ba� ��j8,�+����F�j��f��C6b�ZV5W�۩�#{�r3��L=w�~~o�pk���3+��/"*Ӡ]YJI�z��_^�e��/@Ս���5�F��D?8<QX�ga"��]�;������z.��:_�|�6���X�S>W�;?��{ܘ����n�y��a�s(�b<��H}ұ?OY
���2�!�RwY
�VO���dH�_�)�����R�F�ջw��)��(�x�5�y:�G�L�tՙ�fC����I�����ꮳ��:��t�	�b���`G���g}n�N���L��mh��2c=��Jq>W��M8�WCޕl,<�9���z�*�U7�vm�Y]���6O��{�d��M2�]K���`孫�:���*u⡢�/*���Ho�����;��Wv���,PY_�˖;����J�����k�|�#b�L61��}� ���7/�fI�O���А��1e���\%wD��j"Ma\ԫ�}zeӽ%�,q��8�J�y|_�G��M��V���_u"W2�j?Ҷ~�����2t�(f�A@U�fוK
�"\4�k�U���
�ˌ�Y��Z�z������>�������8�.˧�G���0�t! !�l�`8mѩ��?�½�b}jwL)%d$�/�)���؁���h�\ G]�j/��KN^�6]����W��e�b�r�,��Ҋ����
�Jy�T@�k�����̧�0�/��c�E,I��7�_*����)�sd^����h������;-v�$���{M߅��>�(�~�s�������6�;�6���n�ӧ@�`�/��H���	�w(d�є��ג���Sg���f��z��l���k|���{U�%',yAڐ��a�D@��������7~�ܚ��:|۫6���_�6W9-@WH�+M6k�|lo�_��-'vЙ�hi����9�1\	ө�5��x�5�ٰ��C�A�S!��yj�N_�k�tG^�gM�z���J������ +�C�Q��a������#�g܋���t>������7�s]��_O`i��r� '
q�r�N�2����7�Wı�8��6(�.TX�nV�>�>v,� ��7�O�͛�R��J�h����>s[���6�hT�#�{Z���z2ѝ>.b>7��5Η�����e+ڧ�{�6�`�Ş�5|r�����~{��h� ����v�k��WQ0���N8��;������G���'�ɢ�U=�
���n+��GӒ��"��8YJQ�*�b�Fi�u#�>7����h��\�@�n;:�9!`<J+L���tp�	�S�8A}��U�<�&K�YnQ�׾J�z�}sD[6�C�s]ݣ9y|	�Ӛ���lIô�s;O�Ne�*q��e���4�C��QF(�R��<L���x3��n�Շu?M�q�^k�Q"�Ђy�kGB@SƬy៶R�X��r�϶}�/�X�"]g;4q�C�~��g��Җ��6�s^x$�%����
�:"�^��X�h�.H���ڧ<c�KA�5x�X����H��V��A���\(f�i��>�>
е�m��*��z(t!B��9��9��uLš��CK��N�~YnV��&2�
�^�c
��`M/���<��5���Zu��h�[�p�[!��mA���"XlA6��k���⛧�&pH�(~�S��<��FAr��ťdUH���`�''^�q]~ֺ�Ox�7tɌl���L(�p��v`m�Xu�I�����b0��bE��T�(2R��L=Љ��اns6u����$Q�"�MgGq���N��<u��y"G�&�����9-'Lz�nέ�[���P���`T�8^�0���K�NR3�Xg��P��]�{��\!��X1:ͥ��b�6H;vA���0k�/U�����M
o������S{���O�t��X�� ��=(�o��iގ������ӡ.��|Ą/�p�;3ƕ|{��Y��_��C���dF�{�U�)��y_����������U��` ��;,��2�i{�$�L�}g�ڤ~��BPN3�6rΨΝ*��m��8 �T�Nh�HP�Wi�@�܈,H'���)2K�`u�X%�;_��rǔ̥%����sJ�D}y��-�;A�*�z�Sb`�I�]b즫d�]�J���6�M�����Hn�%�mr��D��r
�ޢ�2o��p�[�	)�ܴ� D��7_���/̷�����v��=��H�\�_���\��2o&K��Tmn�hw���
M�^��</^JH��Q�Eʪ*�|*��PqO�Gq�рs1ނ��F��H�bhsfQ�V�*\���X���5�*�TA�_ˣ��X�`~J�C8�����:��߱�$0.`ʙU�������cڑ{d�� �/��|~���p�oV.�.͖/�S�0PPݚ�ˀ��s�gV��l?���dQo����+ɠ��S���&au`�t��:�iң2:�Z����/-"��4#L3k�_?+��\i܁��G�d��珬����燖�J��f���g������X_+��^T�(��'[?}s����u㎧'50�r�7S���m/��(g	�c���Ϧ��]I&A�e�`S3��(h^��݈c� ��ɋ�a����W2�F�� ��n�B��B�M��K]�xt�r��o)��01<�N�ȤF24%=V�+t-��7�*�١�/_Q�t���_�o�V�л=�!���r��֏0Yj0?Ƴ_V����=2�=���?	e��p�q!2v�q��$���۳F��Z���v�j{��f�O�|��5�R�I/�@�*5)�o{r�f;)�V�j�. #��⭔�I'���X$j��"Kg���Ϫ��������x�+�2S�}�C;i&�p�J{������̅�I�T6�VP��t�c������sm��{�'W<����I�a&�T���z�S��44�L��a�g#�S��\i�8��Ia�`gP�C��Bi������5h?^Ll#P ,��"k��`Oq����(����(A�;١U@����}��~�OX�Х��܆��'�C^�o��QZ)�4�A��8}4�n��䓒��j���p��@S�N:�lm���3(�rM4�V'�SzLR⦁�&H\�Dc�-��b�������Y��>η"��OBT�8Q�t��,�?3���'ID����nhNJpo��L˲*�J-گ�\�%p��~�=Y��!��0v�uh��ǎ,��;:A���s+ۛL2�d���9xK�ٷΘ�Jno���>�c+oA���}9,��v��)hq�/ȫ���0%Y�e����%H����~3���L��c���ұJ.�!Wt�q@�����ܿͿ���L�9j-e���(�>�'L�z�[�"���;���#EZ��y�t�]@�>_нo̯ƶ�f��8Eb����4�����'�ݽ3�ZM���>�3j��M����ޒ>�	!����0;��됳tP<�veE���	�g'I��?c=nGa$XY�L��E���u���-�F�
z�fk*K���{(�+V�Tns�<���J�+����鎸{��Qi6��Zf�=��!�K�\vx���=gc|s#����V����=Qڹ�C��@6��!7{�Ȝ���A�8G�.���ѳ?�2�G��bF�愜tR�qS	��x�1�E]��t��?(�y[����&��������-br�s�>nRCi�/��,�m���o���q�W� `�ܪo�����T�q���>NL�^�\�5�~�W�]o1��v�� ���/o�ϺZ�~�.���l�Q[�)�B�-o�O+X�Hj<�AD;Ez��˝F��!Y�֏����������x	1����K�L�s�m��2p��#yu��9�OOX�U���Ȉ��{���[���>
Ϸ���<�%��
X.���g)�2����"wː�?2�`�V*0�1��	���x��@d�w3� ��Q����8�
��]Az{0��=�M��'Tz'.gr���W"w��{�jR ^@=�18�b���3Ȼ��w��ѻ��;�^�/x*-㶆-��3����]�r`uL�g7����	 �/�`���%�r@���v-��|㔏����Rʎ������HT���K�)��sq����mM6L
�oP�*(W�/C!������������)L9dܡ��l�+�P/�𵫔㽘�Axb�$6��D�`5Hi��
:�Io��`��b�cNe�ll+؏mi֧�r���� �!��}~�@��bO��33(��\(,�z�sW'�d.	�y�^g_�y�����f{��r���H��p�"�w�O�>(�����sH���w��"�]� #����>�2����+okw��07��8I�R��T>��:ˊZ�o�Ǎ^7�$V��֮�1B�l�F (���/��FG!����`�lh�g���=bg�k]4�����F��`�jkW� `��?�D>��	��Z�k���IQ(
ě���QHh��k0�y�Y/e�w�A��%�ӻM�Il����o߬�<�w���?lQ��0���$�>���@ʋQcQ�q�8���'L�����m��%1o=(���c8���?X܄u#x~���8�T�5piX�
O��$~�=�vd�
������\�~@���¹&N���\ԅ$T�O�!i��+�i�Ɨ�3�O�;���1���<��gg�+�,e�M����:Q^�r	c�s�n�`=4��o��k���u���+�ޑ	.��3��� ��Kz�YFʧ�H��T����R�g������4��Cڹ�"e�N���f���S���pO�8���|:e�M��p�R�h�!>S�& (۹�2h6#�hG2
�(�/��˄���&"aӃ��ޒ_U9��8��X�����P�������a�]���z�KIB0�E~�!�7ܤJ��̈l�.���6��z�6���15=��0�17�S�cE�b��K�3�J�[�zk�]K3-o�®�y#ށ��=ƚBu�5(bh"�[?G@������Ppű���DSIAt����z�Fk��<v$�)oN�j�s��m��-��~Vzu������x��e��؇.���S��Q-���o��������j!��l1�睊�u]Jh��*�*D��U"�������$X�R5�7I��ԕ�2�6i�CܲsD[�j�:ʠ��P7����a��R %�xm�%T�Q8��qW�`�)��J]&�++�A���c�E:�7	�i5�I���!���~w4�E�m���� o��BX�@&��KP�h�v$�H>~�#��kbU�j���5�	Y~4_���)K��d8�����d��c��.G��uv1B_�2f����\�W�@��ȌM5�'���Y$n���tܾZ�#d�a�cfy�� �,���T}����υz�2S�X/$�1��d��dr����Ӂ�`I�F��!���#��Qo�����^�A��]Գyr��_��;��
�#:�h��"�o��{��`�>2x�|j.��D�7]�k���D�+��>�9�J��S�C���v�p���c���4=! v���`dN!�3EL�c�J�:�R*�ӌ�?£����m@ۿ��f1��{}y����������8�\��3,~�h6,����^BU8 s���pw����,��@k�D%�af� ?V�_R7F/6��6�Q0?l��ߧK����
O�i�4��9�6�I뼐���k����H9*�*���� U��Z�v$#��S�L��wv�w�nǱ�64�c�_Y��VF}M��~��[jw�����5 �@�0F�ntp���e`���Q%+ �~k�"�)�JAr�d鰔8�"��JbVՙ>{����u-�714���;X����
9�9�I�|�=ou����*���F�4|�3

2��[���AE����AFb'4eD�@�;�����A�k]f�s]tx�.��9R�n�V:,��鮘��\�p���	]ëL`����/!�z?Mx�^��/4���J,��o�xM�yr��V]I�x�L�l�<p!%i$�5P�ɘ��9w���n�j��+g���޸wD0�R��+&�c$r�/�4~H���f���P�LI�*�	���kw�/�/_�'ں^�;X���i����L@�Z���lp��)��>�Rs��∐c	$A���E�1��5��("��pX���rM M!�;4j�\zmZi��r7�΃��7�VA����oB�N�*�;�1QT�ƪV�ܪBص��)^z8~${F<�D4���w����o�=�l*c��Tw��s�.T�<�j�2� ǵ�䕑~ϧ���/X���B�y�#cC E�W���U�Q-ӔS#�(k s��l�[� �L!S���xkq����;3��z�f�IS%�o렭���Sd���T)K2��k_ ������
�Z�1�?>C٨x�e�baY���S5W?Fn��,o�o�W�-i���R ��l����R�ׄM�ӆ:���S���_>Uo�#�l��oh���,='��ڨ��}ڌ%��T��<H�`���in(����ׁ0�osw�d�5��ޘ���)q��7,(�^�t���|��"HA�vz����#&�M�B��d����DB�sȤ�z��z�*�3'V��?�r�ɮ�ґ�
�I�c�%"��~�~�j��{s�)đX(X��Q�$NWk�p%.�t��.�_�����+�Vci��D��@�L-�&L��-��@ل��
��KK�Qʾ�S��׉� ��������V��7��V��0,��{t�-�P\�;�׺��E��p�0�G�=x������D��T�anſG�d����c��I��@�)�붉^ku<�M��
�ê>��D\O�� f�l�IH�׈��V�s�L
���h�+cW��hG��,�\k���̙~�>����'�������W+��@��U��'��KB���ߤr�ߗ��<^�o�[6�e�_�.���}���ڤɉ��\��p_F`�r�0:ؐAF��!aje7�Leg`��>�sU�H!�{�P���C���ؒ��-<'�
�_���s�������"@"̳�"��۞(��Ⱦ�,É1�Q'2%'��S��Z�޺{�Y�������+7��X�h���ݠ	|ɐ��+���6�N��#@zg/�_I��M���
����ɮ�`Y��4o�L�~O�[�^wǩ�ܤ�$=s�ωҙX>`n��F��3A�S����B���7�d;����7�#�7^�z"O����|	!)Q������a}�(�8�"�;:0�9O�{r���Ncܱ�?�M�X�Ý�PaT1���ݬΊ�<���	6u�|�X��+)Dm񟡐5 �����E���)��^'��f���>cPE��A���f���S�Qy��>��m
��Ut���,�tP��S�O�|	�	>�`����A�e����E�N�QR�C�o��lu��\Q"��G"b�B��*��J&�ƨnU�;�P���e&���;�G�T��6'�U�NLK��L�F";_ݧ���7.��6:�����;u�E݁��MP/0w���j�b��gb�ZC�\��+��z]�&y��5��R�ûu��z���h%S*�˛��Nچ�_p���g���V���|���T�I�Nzݵ��"�}h ���o���WJ�Am>_��o�I[�Ӷ��p�q��~�����B����z�� ]�i�'6�3�4Z�����K��-}?�������/6Ou	�Ò]J���K��$ٜ�XR=i����$x2��`�n��-	'h޳�
D'��D��aO�o�b4�[��;7S��￷e�A6?]��ɰ��S�m� -�X�j��BL�@(T�\о�3:ˎ�E��a����e �D������=%f���\j|��~ļ��ŕ�U=1���S�ȍ�:�i�N����w6��z'^�l���Mq����'t��=˵j�n_�צ�]����F]�Y�^}B�p��oJ���!���%J�^�w��Qw�ȧ��G�t�ii�<�Z(�(�_�p�\�v�ȁ���	h�����hsٟ&�/��#܆�cDyV& fI�9	l�ر	a��i�����W��Ee�I[�❩1����T�����qM�_�m�hJq�j������쁽Ǵ��:^����H��cw�ڨR���R�F�+��9�<�ūے�%�����l
�3�� v�ፎb�{�����G�dV|�_�<�/IzzI�q�2��5��|��!Ǯ��٤^��(d4&O�:�hm }�tNe��������Z8�C���\����1ឺ�F!K���01�bgm��.�k�0�\�^��V�r��OM?Pz�An�O>�F��S�}���D�cf�:Œ�O� �O27#��%��P��Q���
��Tٷ�<����:]����eD���M�,Co���^�zL�"p�a�W/P4K<�} �S�Q�I�n?w�$^�Em��#	���8�=��m�S���� V��\��\��&v"x��u�:�#�ij(��_��[s"R��L��D��ǣ����D�`ƫ��X��G���Q�P�0?�S:oNP񺶨�T�z���ڽ����t�y��!ߨ��4Y�v�X��)����$��.�%�����w�ZeL(�9��q���W��T1�y��V����$Nm";�b���� ��\�7C�W.�Vs�I%y�|��X���s��	����$i�4,����haw��3e�m�w^�wmY{b��1\�s÷(3@�h�1�&�k���� �A���7�d��8XIb��Bnwp@*�}Y�{���eJ�id�p��5�/����:T�G���B9�'�r<�f`;��	,���ET��i�6�4�Y 'ʗ��'�3P��5/�3N��E �XK�)	W}l���)3��#"��M���HI�FD��H,�3�fTn �e��!��mE([{1��!Z�Ĥ��)�����M�U⫢�A��C��og�n��(�����rm��=�w��T( ;8	��Z��A�+�ax�6.o~�^����V�q�(�æ�+�*W�g��3J� ��GK"��s����+��"b��Km6R������~���tJ0��|vҬߚG�S'R�S|�Y즴1uA�AK��m�R����D:If�wm5(\�����X����i!7�V�㦯9Y5_�����s?���Vb/nf��Cfs4� ��b!���F��r��B��۽��tz��h������ ǣ:�ͬ*��H�oɥ��Y�!�k3�,�[+��r�q�+˰}8��ٱ�g3�����7�B�PR�ӳ>]����8 ���99~�mRE�y�3j���5�,�j�\��M�$"�� �ځ7�k FBYC�`�^�z���^����}J��X���V&6���aEu�'�R�f�Pa�!K��3��<��Ћ��|z�m��2j`ݷ�A0F^;!�
�� r�K�����V�ف
��!)�5k�#�v�|����Y=�
s���6�#L����Q��#�>���ad���mh������v�RE�#����"����>��+���p�F�/8�@��xT�����OL�Z��E2f|&����pd��,,Ca�� �]���qz�b�Nh������D�ρ;.��u��0Cjν�6�Bz~¢�o}F��)�4���s�A��TL��:�7�Svk3cx~م�N6��%]�~Z��(�=R��6��.3�9)� �~7�V�}6��ioi�������5o��%�S��~Y�&�Lf�G������}\zK
�����xb]"Oy�p3�x�t��`k)%V�Mq��d��U��WP�<�x��<0��㉏�����-��SKT`X�����p����,�����	9�kG\P��8Z���ژ����=F
�m%A�tpY'g�*
��%"�Q���I�B �8��63�ٺ� �~")R'�j�NV̮�M��+��!"��!��3��q?��ݰ���u������R�G'��t�����ؾ�xF���;��`�|&���Œ��U��GN}a0jfß<�%���=�)��0y�ᅻ7�EI����H�qs��('����j��9%P���G�}�sd'���w�/�N�M����k���i������匴��u�s��?f>/�V��"��i³����/�����P��ڤ
��)�AE:����čN3'�AP�l�޻q�+z�f.��ɸ��z������l�#�?i�*~c�����VD�]��m�_չb�҇�Y�����۶�uj'	��LR�o�m}�{Ε��!y��tBA]���-��EG
����?�B
w������߶f���-]�9�o��NB���vȒ��2��ԟmH���69������c[K	��Q7%6%�9�jzNR;��F�:��M>ʃ�o4�}���?��
y�s�2\��<t�R���I�-�L��-�T��1{(;]� P��T ��V�p-�8��j\b\ ݹ�x�l'�mv�A�C[����(8@è�
7]b|����O#+�=ى8����_�����u�qY�D�я:KZ�nQ�&d���>#�Y���"&�1�j,יuV?qr���~"E��x_���"�<��ޘ�yE����ӎ��Ϥ�)9Zr
��G�,���ޕ���R"9��х~���ժ��տf%������%s���[�-w�$�O�V��T�ob���0��-E��8����9������������	�����.����k�H��V��S��д��|�ߎg�y�H��i9SJC�����<�f��y&/�o`m:�]�hK�R�B7E5LQ����Vs�#��C�U׉$����0�������H��3�[�%��t`Օ���.�>��)��\�<~�w߹Mf��wz��!6���ϗ��	Dz�.* 9C;���&���"�+`��Au���.�������ϼ��n�|�8��� =5(�Lc�t��5Q��ڜ���P��NVͩI2���r9�
����#u���0��F�aFQ��-����^Mx�<d�@�g"?}�ם�����B���U����_ � �M��n!�{(���3֫��w[+'�&��G��m���}7[�:�b˸�{����̢�0�����Z��͂��o3(���D<��X�k�(��fp0��MTv���lR��� ��o !9|��*�~�^>�sٿZ�g�o\k��.���e���?�ʀ2 �a���$�eߨ��J����燵2�����i���d�j�ϼ/���S�6ݻ^_$Y��H"�§Bيa���N��(%0�9� d�O&F��r7�����U��9XS���Mg����#XW�9}���aI��}^�8*�kI�m�����CƊ�������ϊP�5A�H�"
|����2jKr�	�r`R�MQ^��eL��T��]��4g.&�,�ri�ӖD����y��/C������ �౫�Fe"���&��K~]&h����AɓA��9�*x���rق.��4я��0m6j�%���{_5��q��OiIw�-�_�	��pkLp$Cṋ"������F�[jj�H8��Y�Y�M
7 륁{��b���s��[��w3��_w�I�Q=�0ű�����k�Lba�#M��0��z�;�$O�����6�N
�%�ne�D�Ng0SB%����Z�:�1�$^����Ddr-�'�	��VV�6D�Kf�0��L[��5��i^O�i����5rj7��<�\��"D&R<����0򡔾�@�����=�@h�Oa�'�Տ�����*N�-����,�����Y!2<�����o��њ�X�Ñ���ח��zp�v�Q�*"
�[?�03@��;l��Y{�+洨���`�ʘ�����!ۘG#Q�9���÷�����&[D����g:�Hn���J}6]�K`R�L$"AbG�-=mo�������s�Y�������;�gi0=�C ^��B�ЙM�Y�\����T���OW�"�c�2eC[��o2)5���Y7��Z��Yx��Ʀ5����Pψ��M�Xr/�]�׶{,t3E�_�3̸�9���e���՘P��+���/�M�Lc�g���`e�o�0��d9ѻ&��h����q��� ����b;�F��D&v����6��Ν4*;&�&Ҥ��p<Ϩ:k���^�!
�¯���������m�v4@FPx��s�<`̶*fS��ƼL"���ŬV����`XC�чŎc6ez~ɏ�9�(�?���s��/7�U�o�Ub�bk*�)����q͓񅬔2Sޅf��A��/+�::u6d�Ao��[W3�I�.Ϡ��j$�1�8$�Lq�E�UrH�L���1A_��Oc��|�
��y B�B�.菕|~�&�K5f�m���c.½s٘��݄*j7|\��$ �������d�l�c���-�FJE����?;�P��P�����LEG����S�kS��꿥�E������az�d.5]�<Ϭ [�Q�r��D����Y��/bTFH�ƥ,ݷ3���QI�8ʍj`@�]�c��=Gy3L�J<��ɘ��f��g�f-Pj-��:M�[�ż������Z�^����ڽ�4�	��Z8��#�R���̲g������q��xe�
���R�fH� Z0��lh���RL�|��{��1^� :@�Fh��j�Ӏ���O��������Gs���1Kf�K]e��������'ȣ�YtvgH�Ft���T�JZݔ5�s���.k]���`����t���㽕��/�0د�s����$�)��,��2��T���Wư�&�[��c�]��/]�dOI8�����4�� �ykK%x[�.�(f�3 B�k�ېX׽�*ZB�L�d*�8o�����q�N�q��R#E�y�P�WiCQ<`|s�\q11���ӥ�����A�qS*L���[��}w"<¦�iCX�U�򷊁��V���%�ʢ5�+���U^-��x2������� �*PZ�'/e6pH&�7�Dt�������faxՍ����PǮ��EBi���)�AqZ�������Yt�@�"��Lͣ�,��]�>�!��<�>
����/�ϝ��3��eb�>B�w3+ni?�7GY�e]#��RZ��4/���<�\D������*mX����2j�%�ϸM29�.I	���=�͞yG.�>J�u�đZh�l�9���-
X�7Y'����b��툨$I����󻓅�8�W&�|^&2�� �bX�S)��X�uD�������,���<�s�VZ#��jA�mOQ�fg�0`�t�j��'y���8X������e����*� F�9���3yU�!}��_�����/fl�Y���x?̻頄F��_���NO�	��M:�>�G"~d5��c�P�|v�8�����#�a�s�=��0���y�R��wE�""vO �ܲE~����;q/�o���p��k�����=��J�=��C�ݾԒ����:�����#ݻ�c%q���4