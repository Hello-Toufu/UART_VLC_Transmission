��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)ND��0Ps�Ke�w"�[���K�g�r�$��˯�{���W:^��jᔋv�#׭M���cY��>f���ˢ�
I�=�����P��:�9.�5�I}�G<�iRI����j$3w����dy\Z"������
@�D������:*�-pw�>>5����y�j�j��������F\.'ʵE��!`0�;K�sq�Cu���Oȕ���j�X=�ˣwXj��Ř,v�E���Xbf������+�O�qy�Ml)1���#u��K�8 xp,��y�i>�ڥ	3��A	�\��� =M��]}����)&���5
���1腽�O��l��<6�&C٭Aь������X�ּs�5���O_zSY^%�2H��t�U?'C����e=�LFE&R$��$�`���m��8�|�R�f��5/�k�#��� p; $D����]�l���Oq����4��o�?��)�^�Ǻ_�CΕߟ���@�k��$$~��l�W�����ju��Z��9���D�)��¦i��?�px���Ƨ�'P�Q���B�ϴy1(E����S���w.]�0�W����M�"�,U;~���g�Ҧ��t>�'8��$8,l��Of�%%u�ǳ�%���F0�
��e���5 �N~B������Z�6Fϙ��\�J��☊���y�Q�ӫDp���f4h�>c��isɆ���%�����wfF�n�d@��ÞR������,���L�Փ:�i��4�H�.�n�U��M�{
����)�*c��"~��1�e{i3ַ�����f�=`jl]0l"2K��j=���q �
S
�����AW;�+���i���j��6B��wʹLHD'H(УGêV�������h�L�z~-ǩ����<I���Z�ȋ6�ºnP�)G!�ُro ]̇��OՏڍ߽��N@S�݀t�-�`��f.,��S��|���uue`�H>P�Td����bOήRZ�I���l�4E�+�2�qLxr7�u��%�A�yKLUk����Z�������r����k�+�4�K��"�*�p/I��q�s�L�Q��&����]�� �7�9ݘ~ʣ�����{4S�拾$���L����m|=SwHT�e̫�IV������o�����؂�X�{�y�����P	����ٜ��!�gL ��X�M	��=��,0��#6�1������~p�NO�#*�0Ƕ!�꿸�T������^������`�G��2�K��BX٦���-'�ۑl���sbӒk�1����x>���#տ��l��
w�[�v��a;<>9�h���������E��r�|~;Vl��-�7�U;��tM��6K�I�{Cu[���"��jj�If��[`�`�hEPr���~����4k�C��&��{���!%�l��C�f���댆�Ŕ��Юu�V�&�� �+�P���	1����mX� �c�TI�U�w��ٴLor�"�85�]����a�����gB�՛�p�<����z�������_�Rv2AΎ~>�Pq�|J7P�ý�/�)�6 �F�1�Δg���=�l�>b�p9�0L�����V*��2�nI g�ՊV!7�(�o�w�ŰIAH�V���Ȗ����ܾT
��֭9���&����i^��JCd�j��xe7�d�Qh��e	�{Ѽ�r�����x	�'}�U�9]y:q��+ ����cn;c�H[��1�A��0<>(n,/����X�1�<7����#��lI�5Ȅ:��ڠ���V�#|�r�>Vo�SϮ�����:^'Ӄ��ae�?%���W>c,��}c�#��[<��F�E*��5=~T���HV�/hD3��Zn���:���*��T�9((#��gU���B���r�f�����0�����)H���ǃ�_a"ڍP���4��d_%?���g߮q�CI\�xg5V��u��ʾM��a������P�9��4m�Vŗ�O�s��8��Av��Uz���Z}�^[M����"+��"+��/.�],�[hU�<�?R��1�jj&p���U5�?����>j��iM�� �C�ѲYw����d���{��kdR4! h�S ֦U�7=ϙM�ґW��ԅ 
ù���ָ���9��'��։n���Lŝ"&"e�t�{Q3�Կ�B�n!�^�����l3�,���HR N���0e�
#ŭMlA(٬3�#
֣��_�M�9[`� t�����\��3���\g;v�*���8�"{}��;~�[p�.�;�W4e��_�ݟ����*JW��|O7GΏ��������o ��5I����Ƞ��������t�oY��h,�Ma%�Y��	�d��Z���Q�ǯt�Gj�NX��k�X�+̼%,�Ԍ{�tk,�	oR�S���ʙB�ǖv�3T���$9H2������3#H�s,���ODm�%�^G|������e�VN��x?aEB�ۛ%+p+�ᘖj$ݭ�>�e��|^���-���j���A�둯9���@I���������A��*ႇ�Y~��J�WtT�?	�
�3��
Ѣ��0�=�<]���}��E��V�ɔ-��t�1���8���FLBP���r74���J��V��ʆ}HPɃ�i!��=+4ɒ�N	E�Ats@�ڟ�E���c�V!}����s90�"������y�w�V��/PvPvVZ]_��\8���!��8.vl¥���U[�RE��@j6	��Rچ�]��_�$�ݕ�!?;Em�Ȏ����?�����IhDa�^!
:��1���(��a4m�s���Ƽ�j	�N��G��/}�_�/C�� Ʋ}|F�D��>�:b1_v[��L���VTE�2Z�� �ґ���67�_�P'�vI��E`��N�F�Ê��o�[�D��
������TmX�.t�Z�������K�����ޞ�%lK�I����}���3��vx,T~v��J�x����o�ZHѦS���r����Nv� �c�7����E��	v�׍K�V,�y�S(�XW3ia������J)�B�f:x�P2�w(Ȏ�W�:gs�ͪh���]��c]�Eo�����e��[c��|��w�0�~n답̨�ͯ�Wu�ρ���J�KmO��FT1P�/����	)�Εa.����	��%I�O���Z�K��P�Sh�>��L ���c�'XnQ�c�{������,B�9�s� �ǵ�n�X�H�r�o:��H���tYw���Tp2,OSC�.��#fS��l�:E��:�W.��I.�Mk�^>y׼��v#�L!�
��<$vz�%�?M�fFG��<���v_�X,#��]#�A�=`�/G�%�oA��@ݞ�<�`� ���ӛc Ģ͂�ܵM���i�|ٿLw�����C���G{�Chq�g2�E��``�`�H��]mX� uWC.m&�e3�H��o}��Q"wE�#�a+����-�L��%V�)����I�jҚ=}s�I_�i���Y�y���%j����*�͞�`�>�J�dW ��k��ǌH�&�t�Q�-�(F`�]�<fX�&�
+�5F��8�U|S�5�-cjIˤ!͉�Ƙo�I��ti����A��t��!�O�L�%��4����sP�L��7_��l�hXYNm���I�ˡ�w�y%��Ħ۲��e�4|��Ҏ�j�LMr���<K�+�轪�J�V�ڐ2�-0�P�p°E[����M,�gꅹ���h�|�5\�ܤ����E�'���h�8��H
�X�hG 3������.6�Qf�����z�=���k�)̰S ��ԃkF,���勠1��;��!C�xL��;V�X����.�¾K�"��TS�M��e�խOϑ,��B&3��Z����t�e��SSg ��t?��TneܓyHJ�f�pî���u+��K0}��oO��H顣v;�Ύ��;A��;�1A �ZU��ڤhkl��fl\�ˉ �ZKx�YF�P��+�]4p�97��\]�Fa�ԣ�<YQ~}Y��94���Jcm��Qc�CC��Y��q�Q;�� �2M+/������Q���jf�ۢ$~���'e��k vb�����~4�я�E`���f7(�6:4��}��� G%��&�X ܕ	���S�x�r;��V���Y(LڼGx-+>���),��q�D�W�_�����L��8?��i�k6wS�:)^��Mà���oܪ�u��7mR��e.l��+(;M7 �EM)�r��a�����W�Q���K�&���a�z]t��ܢ�|v� �Y/(�WDzLT�}��ݏ���F9��w�eW�S�5��z�M#��25S9�&S��$b�&&ሆl��ܤm t��?Z������#�M	��Ҡ�^�=\2�X}����,e�'�
�~a㨕�y���%��۩��}.�o�e�\J�,��Wӈ!d]��q~g:[&:d���3E�K��u�^�	�s2�˛uF`�����J�m$V����PwF�ɘ y���`���Ju	�쨻]h�˽��?M{��`[� ���.\m��W"�~�~0x� {旪�����0�eu��T"�/����z)�RFd�΅�(�L���B\�~��j���o>]ݭg0m�Tb���]�a���;�q;��4������{��U��L�u{�ܫ=�`B�{�>��z=��)eRkC�芥9���ث]cq��r,��\������ݗ��BUh��A�S�}�[[�%u�H�:��avF�LĒ/V���H��(��r2ϼ��)H�GT���7�qK0�`w��Kī�'�ī�Ml�[v�Aq��u3�=#~��R
4�5�i����w��s�u����\#JR� f tCf˗���?H�S��C�R/�Փ�샱Ct�칔z%�S�0?���������=ܥ�y$�Y�M�:�s����t���2w�f�i?�.)o�����\a���D��U���kx.Gs�a��V��~���>|�.��+��z��ZA��Յ�`}�������K�(��N�6�"�'@��ųF����:�qН!���k,X��cE�o�T:aw?&���"О�q�|��F�HZ�!W����B~2�2����<��c�N��6@�n0�� ��y*2��¢7�����XH�a��CD|��fz��ć�ѧ�yӏ�EU�U��Aç){����3�,>��Tُ�����uKP�,�V�����Î�V
����m�͕oM���R#b��nm��}ds�r׹�m@��́H�7k�nIh��di��Wq��EVm�;n�p6�d��m�C~�=��2���S�0���]���r�^��(O�8����4q)�g��|��ڗ����KZ!�@�ALFj�����ݿE�>§	.��`\��ʻq ����2	�5��IP�χ�p��yRIm���y��⺙�q�ڸ*b]�V��y
p1^�T�Ɛ���cz���}���yb����{'�}x�!f����'�L3�Z*y9�v�Ͽ<�9�� ��BO��S}�''�0�����w���/At�0w�O��P�1��ʳ:ٰ-s�S�
�hv��(Oّ�/�^=�;]���UZ�Ѕ�c��?�oXѰ�(�� lq������I�/�ٶ�l�Rˣ���e�1 K�~?J��ia����d"C_�^�e`b.iN��c��u��}K�*`�^�.3^��%�E�����_%7��nX��/�%��[��.}�g�!0H{R�݌~\H�1��Z�'��wLŬ<�ɐ�ġ�kiI�1��C���`=H�I#��u�A��j%�hӺjn�5��� �9iQ8��0�8������Ϸ��*���8"7��"�hf^�{�ĸ��
��k#�I��$Z�b E4f^��s��މ����P4Y�,ҿ�\o�1/�Xz�����pY��'q_��D��.��5��^������NMȬZ+7DَHRq�Pe97�8?U�������=7x5�M��]$"�8zv"�+�U�;��[�]cm+f�?v_�m��DD�V)	�0��GH���z����T�q��-]�f�f:թ��pH��č�s�s�`۶:e���T$[`�io�srNe���cLT>�sۨ|� v���H	Vs̢��[fR���h�B�v�_���*��}��hmN68\��v4�g�$���8H o�>�
y��۟s��8��U��.��/x)���g�"M�� -o�+��ʂ���`Ê���\�H���,s&gQ*=��W�C<���.��MC (��u���Bu��U�8A����D��-�_�t�ɮ@L�?Ȱ�Czk����(8�_FI�Rr�H��m!��k�}��G���FY|d}�eN#n���*�HN)T�>���������i