��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�G��ˊ�Q�+���6�k�̷mX��7��]��Y��F��1�Zo�F{��F��$#	6G��%�Pi=��'&�b4*) �v{1g�'�}�(���G�A}�	�:��Dn�V�Gܶ��E��y'���`�3%B�Lڎ�*�-��kq}�b�q����5�\r���R����IQhie��Qj��G�Za�	��b"Z���Q$�Iuw%HŢ��_�F �Γa����i@!�
��@ w�i9~8z�,E�ɶ7�;���T��]Z��X��¯]΁�����~�V��}�E��8��R���B0ߒ�:��ݥ3��MCM����x�#��_U����Vp��V�j����>3:�����bsa��i��C�ܨl%�zQ9Ü��B��%s���[&� ��K�_9%Y{3c5C�Ju�+���;x!-%�( M��*oIv�U�ŭ6F��,P6���l�{�ҧ��J����*B��<��R���+Z;����4����a{�L*8N�K~��h�y�Iq�F� O���6�eނv��I���NgCY
�ހM�6v�PT�k�;�4���,�YI`p`��eT�q�p`����뱘UP�|��Rtk�w�1aڼo��y��^���^�P%���F���p�e)V)�.��{�G��fZRp�'� X�1MT��WY�}%{ᵹTu/:�� �1\��W#��C"Ph��`�����2`����ۣ�Y�v!��(�+,�e��l�K/2�_���]<|Nv�>l ��0{IRt1P3�I���7�v�;ش �쾲��=����}����~���&1�
�%y��ZX��ԇ99Yx��޻y M�*���gL�����>>6Q��&�*��X%sX��R�=�)k��~�Q5<�DTS{�d(�n�T��nZ�9����~b+���o2ɸO��)�O͓s@�V�h|��N�߻(]�Y.YZ��
����������J�ւ��b
 '�Ld�{T6���Q��A�˹�p����Պ�����Rd�̖vܷ�9f\_--�O[�����m�7.�5�W�f���tZ��<W>y�2ag-�@:��^���F�`�#G__����ϼZ.-<ηǻ�?��Jh[����*�XA�ͻ/h!�⠊��V(d�����g�����_�.�$����u����F����˕�#�"=kalZ��8�Ye:�k������5=4@gMH�i~j�0�w����WI��d��I����<���dI !fg�Rݬ������{���y����w��-�s � �kG�rb���% �� "n�-Kφg�5'bu��O�3�Wq[���*�F�X^��w���B���O��kS%��l���<����Дę`�O��z�$�K�t7ȿ��B�"F*� Մ_�xkZHӱ��+ �/7���?�/f���y_��u'��|�J��D`9v �}:b�4�ƀ�p��i��F�ʟ���Mhy�	&�����: ���e<F��
ҫPM�������n���Y��[��I6i;�k�Y]"~���!��:�x	�6�*H	IT�T�9.`��bWQZ��M� �sq��{���'R�Ow�*D[�2���Į�S[-���YYi���aU��|��uA}���y���}�N�s�V����[�5��Y��ֻc�}�鱁����L0�p���1�;d\Q�ؾ��b7p:۵��!)�����bA,f���&�3�@N�ߊ�.S����i��^��-$x���%��b�$~7��X~v9����,�O!� r�ʵ���"��oC���F�Ƣ����[TZT1�ګ��β�Ѷ�ݮ�w�y�j�X�n����f�Z����'=G�쟲d���
�4�Ҷ|���Rc������}�����gő������Be�� Pv&"�X����N?v��H\[�x��U�8� �ྐྵ�[���ӌʁ���-	հ�eƓ�����9�p	���X�ڇgh19L-8��Z�R9>�ئ�&(w]�TV��X��%�mw8�d\��f\����Ȅ7;�λ����Ԍ�2�[#�:j>�X
d#oJ�(�"�l.)����,6�
��������Ur� �^%��E��O$ibNy��N�'&��?>;O���3���=�)�:P,]��Sa�s��<�`�_�i������Ɠ�Ef�������� _D��ܔߨ<�(Z�̼>�J%�!�>q��`�-ϩ� ����kt]��X���<��!��@��p��g۪�f�?1ۧL�o��t���*=�k@B?��e����b8�ͧ��$�z'��٢!'�E��j�֦�!�F�aާd'g�f	f%��5�sФ0>���3�chiMA}�cyC�	�����qdjd��>S�]���9��xLw ���E0�Z�q�*L�D�3}���q+����v���=h/����$�Q��c�x�����T�@�1�Uf
��ot;C�r�8���^C0� Y�1i-^�l��x3K�Ԝ�;���O4ޙ߿f�R�1)lڡ*��m�;��E��(Ņ��A�Gm�
F7�'䔡 �Iv��4����k+Lڕ>3��*7�M��P�2f��>ξ���uR��&�	`"ݩF�,G�B��UmG��Y`q!��E+��F]�P�R$B��ܘ��'�%)�Kd jp�En$s�d��B�5F�s��V�X��)�rú�ld�չ��[>�����c��`����, 66 [r��I� H�O�j�69�;���bn���+F�H��r}6~ۦPQW���%��((��]�?�f�\K�ć��=�}�ެ�L����i��B7����W;��ʲ3�W0�7SR���c��X�N�������]�nb���n�(��q�Z��/R+����q*�����[$�rju?�����m�V�S�y��P�L�|늶��?ѽ�G%V� Yj�C�8� �ir��Q���Zs�4"ү����#5��G���>�n��ƭs����8a#�����g6~�6��w*�.��w�_�2:۱��:�~�M\�>� �1_[ec捪񊒑�Ӎr�i�\�����7�(�?%���/ԨN~��r��?��B^��&K|h���(�i��#���x��g�����
9D:�G�⫵��/$\�\���H�C�M��F}Xj⦁v ��7A����)��b9�k�ԫoynt���k�""̛Z���?�U<(��q��p�I�ު�(|��wdST�rv����3�[a�8�k> :8��?A+�tc�|$���G�r�g��xZ�<]+E�㬗��ۡ3�Y�!`CJ�IS�,��ʨe�&y�R�;�b��9�i�D�~��Y���hd��!���.6�j�+Jh���׈��K�k��+��0���v&�(�����Fh˞�|kbQ7TΑ���b��%K �H8�Cm�i�)7�xt~���ü�W��y@����C�� Č�7-�����8�_cblH�
s{��1����rd��_��8�+�ʝD�>�	� �2W�,���G��q7�R�۵w*Xb�k)Kbed��M����P�K��B�Ff�?�XQŖ���5wb�L�G��"�?I�~�w������ڃZ9
%�)�ƔAWP��m�E���	�@hF4G@GIw�`�U���9^�=%�eC0�}�a\�ad)m�k��FSs�c&ē`����GӘh���X�g��i��]���PГw8:X�r(�BZ��4'�60������(&�8ap�CUL�};$%>��������^?|0Xf��\j�����?pr���*�^G$����w��[x�F�`��wPT.���6���"n!��`�m�ay��c�T.�0��������7�2�@{-O�*f����f
�ea���K�9�Z�g=�K_X���'����Q��j�C��^߳]���Ψ?s�3���2+���ìH��Bv��+v^�R^�sG��D�X�@����@!�h��(�6e�D��F9�l���8c?�B���ޥ�$��?��Dng�ur�e\�2����c���i�	`�Gq.����ӣ䑨�T@���]�fy�	�Jl��()��`&k�T_���i�j=���o�{�Ͳ4^��qG�B)i�$J�u��~�(�ȆO�"&��L�u�:�%�(?M�)��%F�L��q�!��cn��j�qj��%:��&�a�T
�j{�:Afa�4��f�׹	�LE,���3d�����z4��;v�b�]�wj,Ʃ�A%M���@±��<:7�2����i h�HQp��G`����C0��
�"R�+���ިH��XgK������Q��r4(� ���L *�8R,��D�聱����#�}�Ӥ�00�፽���u�/�N�3���@8*�.s!	���`����+C�t��Js�(�Y�oY�-�����@/l�5k:�%��d(�������T�Þ7HKJ��Md�:�T,~���7�= Ie;��jou������֪���~�k�=�I���.�a�~"ˆ�c�PR��1i�X��`k���Z4s�5x�2�|L~��e��dؘHqA7��SS4D��L���t���M���	2�!&ͱ�=���g۫e��"�Q�Am�~�t@�2q�s�Bk��.Î�Xp�|� ���԰C�UJ�p
�q�%4��L���p��_�jV����Yt+���>�
��UvI���8���q7H�-*��D>'�9K_?�Ow���G���� \sJm���{aw"#�d@�R�ݹ�"�&��At�r�k �P~�`�'xJ?<���9Y���78ۄ<�+�g�[�nw�t`j�����8��:�=W�����g��*�y��6��ӌ��D��.f�ד�#m�,�M��Z����ǣ`Ky6;	ܴ�ɷ��� !����D^��,�RS�3&���=ĔF*���c AS7�ê]%�I�&F5]���Em ����·gRf$7g�;} �3L��B����7�f
�� �LJ��K��=���XLqU�����+c�M�S����;\��b3��2��)_���,G�X~&�G(� �´������J1.��a�Tg;lP�OM��p8K g�I2�xno89[U�\�n��Wr;Lt�,��M�����I�������2	)�H�G�|K�f`���К˲/'�Y�t1��AqK��`t0lXF*����
��o˪���]BO*�ɾy},�DGL�w�E;1����|=��.���1��U�T۔r��hV&GT$�, �ќ�!�5ȉ{�M�nRzK��LqGV^P���������MNZ|��n���q�[���(��45����M��+�w�e�!ِ�,Z��S_�5]g������-�E S��8`�)�֭�~��}�n��ѯK�?�bx2kN�ZHV4{�e�%�ӛs���9�$���������Vܱ���<UN�$cJA��u��<�����L��B�3|܅ ����я��o��OaW������0��������D����%��}UE"@�z��)bW37��
��Ee\6�������s�8tl�(�?Nr�~�T�Ǟ7v��I1��S����ɭ��QD�h�8��S�1��O�_�?���/��u����t|r^V^�Y�$AL���R��1����S9^ݞ.[5_��߂a�8'�a�z���>J�C���6�x��[D*ki���'�U�o��GN�&�F�lK���������p`itfdk%?p1z\��h�����&���?��)�&�	�H�y5"�.��o`���UW��&7��?��9I`ٹ	����^�ܷg��u&���M ҤF��O�R�r�wJ���S
J jq&�Ǣ8#(���y�Y7�����1z�b����`�%/�38m��7nЦ� ���+�o�D�����wo���K�ͩ5��e���C;9$sH�)~Px*�(S��OM�jB�b^����)^7���d�E�Uz������8�����nQ~�/��"K�	@w~Mq{�ȸB_8�PX_������vq�U`U���X����r}��S�N�zHT���e� ��.(����k�/d�*#ӛ�u��n��N��ц�oI��_\>�[/�Q�mp�Mˋ���Ɲ!ށ��sS�4��Ϸ�x(�ң�E#<lN�^\�#2�Y�^�;����+(S8��)���РGs�1DA������QpG��Q쯶3�b��yn�T-;�T~V�9��K֔����ԝe�q�(O%+����}H0e;�j��;���f�KO�3P�)�k�0C��F����I�o��B�����������Ko������}�p����z�
����u_yBl����?kS�sޝ�:B�G�Nu�:��1-*=�:%��[�V���!���A�q��p�� �;kK��q��ɁR���-,���#H!~>�}���ᨙM0@�T�v �
)��=5-�{aYSO����쎷��v7���"u2�э�4+;�����u)q��h��_� ?N�>�*G�4B�����Дa:�bd>�`$�`�VR���@c����@�a�c��I!��hM��H5.�]�ԼAh�; ��N����$ưl��ɥ��~��1V�P���� =����נ�d�h���z�K�\�~7�|�h|�vr�7t7�R�Y���8oEYvȕߥ4i�V�w���b��k���9*�̙�;��ϰ+u�"���"#^�����'1-u0
�Q_�¹�:R�v�K�����]
���a��a��T(��(]������w��a�z]�6�}$�X��"��}z��>c^������u�?�������z��Y\�e�*�Xc�dbW� ~	y�A_!�SGU�E(��(����H��eU͙�6s��a�p���Z�Es4\����9�� ��,����x�fY�Sl{��FC�c��@��-���;8\Y��I�C��(��󻸏��'��LM����w�;�̌�e,�]ߛ����[� ������?��Vt�l�E�qx���K5}$16��x�7>���G�vx������о|p����MBU|�ֶ̾��ҳ��փ�q�#�m>�0�F�B�w�EIنsu������Z��DL祾���e!S��}k\���7Ж��f参��!b���ˮs����x�w;)�a���U��Y��0={������Ҝ�J��1Xwb��[�j�@]��Pz��k_�F��Bأ��e�o� =+���n�Tr*��+Q{�i����gSڙ�;�8�a�>E�[ ��B0��6�u��3ixW�_�R���H��3�2��L]V��� 6*N�KS"����rBX���g��K��A�[oZW�-���K#����-�����a1���N�M�<���$�����+�y��Յ���kz��!%�<X�1�ɏ�삑V�^��=�gg�}.�I���tq�.���F��!`�8R���7�l��]i���(ˁ�H��������gyl���&���J��[h�X+Z�ش�6�j�Q�՛��e���&NN=/#y4�����3]G;�R��,�+�X�-���C��M�<e��l��`�6E�#�tTi_��{�g�"�7XD��'9��]�<`?y��նP�5fz�lS���v��v��e��XG}N����pRNK[����`8)�h-F(��:ͬ��aMܲMR����:o������G�7������	�/VׄVu�\�45!�I�oyRA�Z�����Fuz�g�R����{��A�}�9�7������^�:d��]#�F}�÷��Huv=0M�����wq�%\�\��;DP����1���g���5E}��;��W��j�I:ӽlc�{?�X�:�yirxY�����
�FȲ!uv�	���w��Hj�,�cը�̍�p34���&ڡ�j�d�!<�`���߿�:�'W�p�h��`�_aP൝>P��@���Dח:��6�z)�s�sN���;Kn�|B��2�ǬŜ�9evll���W�%�I�]
�@;06�pΙDtB��iCj�#�[�r�)��x��8�&������|>a�F���	��akw�����I�{�:J�ə�����bGV�!J�0y���8�d)8�����=����h4b�W�ATL
c]���U�_y��k��Ʌ�l&Aי�LmZ���Q;&E%���?�ɘ������ɶ�NO6�p���[�H�7��n�����aC���I	�J��2D�K��I[\�4�Xךa�]�U��
���.���_�ӄ,�aGD�^�F�Gw�(3c���W"d�T�ƪ�$*ˇ><R��72�݊���%#�pE~2�[���ī��v��+~\
5��F��Fg۴�Ôܘ;�^΢h��ַ���.�9c�rvX�R�����r��{���-��Q(3M�v�^TK؟�:]���&�d"������@@�U����gq5]<7
�� \I`\�����
�Ա��;�^�YK���b���:��ԂyM���Ȩ� �`���aJ����z��ՙ_l02k���_�הГՖ<c���{9�� ���#�:)�6�3P�z�s�~t
�2�0Ι���qJ&u�j�$v�l���Xc�d���ĸ�.@-��s�0�e�"v��4.؇��%=tj�u����tZ��C{[������*2�j�@Y�Q�_�� �U�Ie ��,e ��d!�|�u��Q�fnUP~0� ��uc� �L�b+�3$���� �-�j��)3��XNE�]�,�A�m%�{�Z�.��N$;����M}���"�X�	�C� Ȏ��d�`g��^/�Yr+h�����ιtK�pش��h�O1�f�=샐�l�1��cO����n!�|�F�@a���£������b��t�J}n�m�D��^,[)	LY���x$ k:��p���
:)W8���e��c&�wf�Ԛp7���a� �o�NV5�ܡ3ĳL��	�=�f~�ɫ|�Ds���Z��"�2-~�����"�����d��k�I��n�+��j�凳T4���l�-qc�0\tҵ��c���w���� �\��;4`��,}���I�ڍ+�9�\;��f8��$�~Փ����i ��*W(9�*e�%
A��9w�3Ľֿؖ݊�ƶ_�������d��ӈ�g��**��)�������'ag*�r��fUV&��Y�r������1��)U"}��4�x�@eRuf-�F}&\��Q�U���s��0�] �ϫ��?�i5�{@��֙b_M�8�5�1>t�Nz>�&��ۑDo�\!�0r�G�mRǳڗ@n	������e(��lt_��衸�@'�� ���Bxsޑ�����L'���M�s��.�0����I�L�`���K��4�C!-�۹��k���Ϻ��>�_&���{=�=�\�)�Y�,8�H���Kp쬖��<cΩ��1��Z���-AF	��<��������ڍWV�t2Ϣ����*�;���Ȝ��}���/���y[�=�sP4UٰI-^T"�j�}�mDIQ$dC��y���orj�N���|��|�ADټ+tZ�J��0N@�4R�tzC=ꀫ�?��O}u��*�Ph��{as��F/��ޤ�xf��V@�PXv�}����2��Z�%�V"Z��Ε"�2�.x�8�Y�{�;�=搩?��;;z����׶n���1R��Q�=�:άH��i�J�!�o�[���y'W_Ǻ]�RkE�{�$��G�4��f���h�Bk-���#O܈�ƞ�s���<�JO���?�͉T��?�ھB^�幄(
� Z�l컆㪩���d�D}rv�����W��sW�4�z�O��pΣ���)���J�ˢ-��t�?��}��'���d0���Ex�����%�.����1Ś���$c��:��C/�m��u%4��\l�1�Esﺈ�ͼbS��K��a��ò������f��y��Թ`_��f���uc|떀me�wJ3�