// wait_time_threshold.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module wait_time_threshold (
		output wire [7:0] source  // sources.source
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (0),
		.source_width            (8),
		.source_initial_value    ("40"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (source), // sources.source
		.source_ena (1'b1)    // (terminated)
	);

endmodule
