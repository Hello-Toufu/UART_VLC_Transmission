
module manual_rst (
	source);	

	output	[3:0]	source;
endmodule
