��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)NCA���ɠ�?� �Žw	�h5����(Y�_t��'�o#��6���:�i;a�*��MO�[�&v>z��?2E0e�U�a����W|Bӹ���8�iQ(wx�?��*]KS���T�7vw����dF)eMȥ���|���I��^����B������0�d�R0��f/�B`(�[?�\y�,l7/��,.%B�!߹�L�]�B]��=�Aؘ�ÙVzJ.�k�=�4x�Mh_X�ԯ����zM�F�R�R����2�
%ݱm�"�X�K:��� �L�������C�_�~�,��E��J�w=KA�1�0�8g�_[�4��L��Y���A���0f��y-�-�1[Ղ
h���ɘ�&/��9��[I�
3�!��6����*������u&��O���(gwʧ���`�1��/~gI���;�>;�D�O�ɀ}�fJ���^w����,��̮p�N|���N7ae?F������T۸�H�M��ޒ�ǝ���i��*�nkVI��G�M�a�dQH%�EP��J,����lcl	�~>�c}���ߠ�)�'S�����5|�&E�����+�c� `6�g���XW�F��	�#\�P?�蜋>W�l;"�r�������Q�]�eU��C�ڝ*��'�㶇���Ď# �obJ��8u��&�{�`�x]�^&����x�.��T�,�[Cr!�T��9�3�VI;  ���m��|~�8�n��p��Ғ2����֜��t>M��m���r�p̾?\A����*^��`� س,�"���%a����)��	6o���υL��a�����7�y0�0�sP����;��ȴ:[�jl b��m�Ws0��Xz2�?���0z�թ{���8�N�T-V֎�mL���$��Ͻ�����.�\���8iH�>*�����}�7��D��߄	���#~���بW��ϡ$����}]��9�K�"������}�b�43^�oE��,o+�+ac��1]e�A2X�/�1�59�A��6�^ r��¦/(�)�HR/;U|Iв��i^�;�+16O{Z��txj$��_��_�ՏF"�Y2��(^�c�����[�&C?���gfɢ��{�����
����g��:*����_��8�1=)q��>$n�|Si$	�8���k��(E:���r�L�$�}����_o/��M��TG�'�j���P̈(*�dh�$�ٳ�N04��= �*`>d}�'��l�M��X��r:����$��S�J�{��k������)Ap�v����j�e�����?��FZ�-Y�F_r�>�5���탏w��*����ᛙW�s�eo���`�-���\0��������?�%��u
�����F����	��{�S'ҍ����i�=��jM���5�31	�Y`�a"B�,�\����Q�]�����~T��������qVC2펅���
	�ݮ��I8�t�UOdŹ@����$|�u�����	�_�<�~�6�s�FS��y�`��\o+��s�e�l�2�t1Tz$b�(�s�Dj'�S�
����A�+�Ά_SƦ������͢FU_ŵe�Z/Q��Ă�V n):P+�Nh�Q�P�*}Y��g�Zl?��0Ն�"�$��	=m憨f�����(��4q	?����B��^�1�х���k������܊K��U��tG�]4J/R������ug:��������=��M��x�n����U�&����~X��!��LE�����V�����jf�ݣfn ��K��gf�D�*u%��]C�