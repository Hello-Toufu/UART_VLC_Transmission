
module wait_time_threshold (
	source);	

	output	[7:0]	source;
endmodule
