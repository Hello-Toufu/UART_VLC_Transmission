��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N'�|Z_&i������w�M
U*C�����H���t#g4�od�D*2�}V���F����9�an���+U������Z����7�o�&K�D�%��t�_m�"89���km�[��<L^�� �l�3=Bh�A@�\�#=蓝��Pk��L:��|�a�PGjV�5Ow�Z�jd�)!$�ec�%���Y�ٵ�T���0�϶N�B�T��9�b�4�?H���ߚ�e=��K�, :o��^&S3 [~]�~b¿K�A�I�89
Mr,�	�U�)����S��R�#͏I��@y4
!�w@!�+	�Q�Խ�����t�=c��q�g���	��ZH�3?��R*�(�D3��n�_���I�C�&$]�ߔ��I���!x�H�����9>	��S�����Y(�$�,Iծ��ȏD�T���J��	2�0�M�P�>x����Z��Q�W�o�3b�6�� #�޿�I�'߿�_.h����S<�Nz�>���/v'�_G"ʥ��CH�P?/΀	/ �+�����9mW�����������c%�A�ٍg��G���g��S�]81G>�h��x�!��c^��"�7�ä�b,0��CT�����u�������]���_�,��u�u���k	��klQ��G�:
�������`m�{|\�߬���
?�$a��J���E��:6]��PӝJy��:T��0��(�ƇUy���Z�)�e�8��!J.o^$<��{�H:��q�����C����_�����7�v��*Y�w�����,0,�����e�۵��ݷ��X�0Q�@������<�^�m]̈5]�wR���#���Nm�����I���J��f'P�-�@[p"K董�-�n�tR��K��@
�K<�|�y�p� US�\p�vʟ��1���.S]�D���{,��5M:�����im��pC������Y9!yg&c�<#BQ�R�W��N����Pϒ�]��P�_�V��v�P~0��?dJկ$��j֝ ��q��!4��������r�������G��$X�G3u�`,ռ�A��wǻ����j����OT��!�Ŕd�5�3tѰ�uoLuц=�����'� ����t�H�����H���������'D��4��+��&-��u'EF����7�u��a��6\�+�`��t0ӡK�©3S�{+)y~�U,OܹgD���j�:�f�/���Ҩ}��=nW�s������ԟ:Ǥ+����q�2�؃�H����u��Ox�K
�S������8@�7^h#a�P���nO�4�%�,<o���D�:`��Y\ˎPPM�LXl��~�~c�mZ���X����ʮ�m;0ס��c^�@��ө�O������_�y�P۹�I��ک�-ު�3}�ce��&������æ�0D��4�e�>#'�������jf9�YO�2:a2�'xP'8�
����Z꿝3B)OXҋe�����a[mNa�����S��c˅>+�<_���m��Q�f�^��mED�b�{;��!��(Zĉ���l�H����B}ݒƮ��b�FT���[D>��	�bSI�՗�Pu+���C��l/2 �W�3h���{\k	��s�L��g5S�E�J�?0h�E��>����9R�Yq�YR.m��2����Xke{l�U�V��ܯ��� bs���n�LGx�7>A��;��U��y�R��[����0]�xJa4����,,�e��89�Ej@�3aj:��^M'�t���$�vu�W�߬����/���Cӵ��^��Z�s=�`RxE+�a��
�Gs&㦴�v�:�ꫪGR!�8��8+��U�Sc��^Zr��i-�q�Ӗ�S��O$�A�R�9򙔯 W4��b��8N.��������K~�D��0{���]��P�㢍r�Ҡ�f���D��<��ll���_T�AB�X�{��(K�W�|�7� ���R�n1%�z��z��w@%sm>B�,�#|�K�����V=)tM��5�ȿ�,|_����`�)��~eƦh�����p���MO��V/�G�×�k�.�5�_Ԉ��t/��K��?�献!�^��S��XK�I��2��-������ӌj3BU2��A��e5M)��~�6=/R:J^F�h Q��`������y��.�A�����Yomf�C�g�VYW� ��#�c#�2���\�p@b<T�Ͱ�4��
�^E�m�ח�}J�/Y��Z	
�H(A�&�~��N�������d�)�Fu�']z��*�V���_Mw��}�J9�3z�ی���"��(�z���$lC�bh������Y��$RC@7��~4cˌ2	��}���`��6�(3��Yn{�RD�p����$�5hVZ���
�����m{̯�¯�Ae��RѲ��DuX������^�	�؇���^p���{5��<�R�~e����>��hG�pS
cj��_X$���	���,"�uE��J6�:eU��rd<����%����M�xR��g�7+�'Bכ������)�1$W��<������Jz�"p�����Xeε6lvÜ5?�d�����D�l��W,�j�ߧ|X@���5��?:��.N�Z�Ͼ�"����b��B��yB�.�b��u;���ɶ=�Ğ��ϙ(����������Dp��T�4$*��WG�S�U��Ag��>��QF�N\U�b$���F1͟��h�蛁�Lt��;W�A4Ui����*W�h��XfƦ�<ԛnլ��K��giN(�vR�Ӓb�<c42�}���ĵz�E�v����[��rNՐ@�ZTX��FO�k��6���iM)��	��nKVwuR�$W���(Yc�*2Uc��\Q���C�*)��Fˀy6������;M�V����YT7�Ny�3`���NYW��9����6����aK9�
}��5�8��m�u���@����ʹ{}�Z���S�M`Q�{(DS��s��'6H#�˃��($ppC3�Ǹ����Q(�Ρ�;&8ΉN� �*A�5(��(~���5�����J��Z�F��ڴgh�7]ͮ�w$jI����+�����*_�K_n���`�L�Cs���9�F��������;xsgM�KN���^ʑ4[��;#z�� �{�����z��!�x�2�%l^�p��9��׷''��kԽhUļ}2�8�9H/�Im)j�S�<z�U�.H�6�:�2V�1τ�e�Y'�s����r��١����^ �n=�#�0^��=3��#��"J�
H4&C8��a
폦P$�$ؓ�B�/�}�k��lZ����dD߀��p�B
+�n�k�g&=(�㪅��U��I�c�<�/��-$'��!Ng�_fZ�'���w���KzD����9�s)�2X��Z�\)ӌ�%��+����~�/�Jl�QT��c�gqx�n���B707e��t��Þ�~ǜ=��5�$�d�5*��o1a���y��DvF92��Xc��E_~ӂx�^����g��@F6=�$�C�C������L �����R�╧��
��0�oD�,2�i�)��2���p�{n��W�4�{&�P��A�\�IK�`��`]�L�3w�p��FHt�DNDEg�37��as�K����W��tǷ8�®8��w#��p3�'�ƪW6�����RC*xEr�����dhG`�W�Q\:�����s�o�9��SY����5^1��m��\ny�l��ɖش�	�q��8[
H�ܳ6�7��-���3!#ʶ����_"����Pk)&�yab����2`�o9��&�M�b��~�$Uv��,��K���K�����Fb�k�k��.څ���1�r���H��SQ��~�{$����<1RX,>�uv$Zo-� $�9;R 馰�ԉ�͵Qr�6��Ϯ�UӾ�p��2�Z3[h�����yi�\3��� ��3�vE1��ڱu/I����G�A��'�r�@�K�(y@"k(����Y.��I�!�׏��z-F,�s�[f�!)�O����cS"kq��x�x@.�|I�4�\�AyC��2#�Ŧ���]h|g��k� �|%DCp�i�K k"e�t�ѧ����7�?��hDT)�Z[�a�em!�팭���ax��c�j3�I�����<��_'��M�'-�����ۃ;F�fQ���~��B^��QO�v
��MC��`���`3�+A��tB/��u��!�{�wZ례����]kOB���ZҶ�?g�&.�����f��BV�?|�o���J����a ���P��6�s�ҿ�u!��M�����dq�+oa�l}��|S���Hx���J/A�~�18������<\ׅ=FaI�ZJ93��Ym,&��	jlp��)}�&܆��/섖(ϼ��PTd�@���������<�� �ۚ���-���D#��>ٲQ�,e��&^ǥ����H���2 Ĉ�|>�N²��<��/[[���M����$�)�N*?�A����>�J��{L�,���4:��7�N �n�Mx,շ���+k���o$����Zb�T���`��t��u�z_a�d���a�|�O��O
3/(ZJ��%)+m3+Z�I����t�
tF�����i��%W��ꕐ����],�k�O��Q߭�p���z�S��y��E�����y�&�qvD�K�<�3y�;��2C���^���(��h{��Rp��1�H�����K"SidO��Q��,!#����}1������w�a�k����G`�à�z��)"�T�X Q���3�����a<��0�̝�9D�p��X'z���l�j�F��������+��y��t�q�J1�Sq�&g��A�R�H���ۯ���5��0��)�IkGH��aaCwYܴ4�Q�l��:��җn��1����5T��.��UӾJ y��+
nZ�k>\HvA�Ƕ,�X�'pOjK������NpH��2����ҫ}1J�P����*Vi�q�I�$�8�0v��� ]�M�b����{	^�����0��2n�/��^��D�"%&P��6<.|D�_��5D�p�ʫ������+�@�&�&7u�tX�أ�υUx�  ��S���y7`�e�ڷ�p��#�ac��	�XҘ̮�5 �2�!:��Ȅx��N�r�B"y5-���.�fR�� �t�4�-�CȽ�8a���vy�(��+�-Cׯ�����(�gf��b�DBa���QD���Y,	��b���:D(L���:Ӣ����y.t1��$��*1dQoE��K_��#�B[�a>��H�Sl���μ)��ֆ_�A�
Ҋ	��`�6��ָ8�sasg��Zv@�0BO8��n�V8��4�-
����V:����sP{p^�&�����������X)]�P<*�G���j��m��M<��E;,ūc6�W����tZ��"x�M�H��հ�j��kvmoKl�� �Nbil^�1���S�&���sd�X�fC�F��"�ָt���1��g^6��Zն0f�W��.����\�PmV���������ڬ�]�>���	�i�|��B��(�23����9J
 �ش��:���Np�
���4 2kެ:����_y����.�Y*�����	.���\��!K���K�A����H�V9�����4oW'G�i�~2���0ä�5P�n�Y�0[�z�J�F�?��T�*gA�]qs�&Ox���\�n�dc1UM�PI	��l���/hZL�d�j0ƾ<�L�k$
rgG/R�x��b���\Rj.��B� ��ѥpoo4���L;�v��74�'�A,��0�5�X@��?����pb�#�^m; !�G'��1�b���Xng/%�g��ef�XYʠ���+�`-�6p�:�Ѧ' ����3����G(�?U�x����v)wYȈ���ʱ��~ţ����mF�.mu������-Ǐ�8�'�H�X��������eu!:s|�P4;f`��N���e/#x"���4��iR��G����B��hl��u������d�~��rN�Ȟ�P�WK
.���	Gvh���ܸWt���������\f�<�J��kQ������o.6GE�}����ש�f:��@�����[或�/=���>o��``�՘F���ܥ�k"V*�\4��P`%F=PsFfX��I�=��CT�p���~:������Rp�^1�}���,��]�n�/�� ,H5���.�)�pSZ�U�$���XC�[5�p����=�-��5E�䟖b9Ҫ�㨹�G�C�L�j2,�_�,�e�@�+��� �;_1�qEm��-D2�Ku��̭1���z�P\T����u4����� ��Q��h1O�'t���`W�U}+:�W�Ʈu�
ּCżA��L=��k}+�J�W����%��d{��D7[(&̲��HcI�p�D"n��$?�<�3d�_��:�!7�G8��W��7���<���a
|j��ڨ �jۈp���j�ƴ�z� ��s��a��kA����ŗ4<v��-��U����Es�jழ��{Y;����V�K��"��h	^�n(�R���ĊB��QmH!�J0���K�9	���t���2e:�`*M�BzᠰA�ل��3�lZ�=)����K^)��Z�H��`���"�����~<��ej��p;�~#����a���̗���	�x] ��U^r@n��&����;�, ��Ko��U��jO��]�oLs4���ĥE��wE~�Q����ɇ*�H�ȆSM��4v���Ȱ贱�!?Ja(M$5���&�-��l�[�`{�3(��WHް�>��@��jR�$�l��ڭtc�⹼_��J &���5������`��D�ڊ����pM�t+��#��h�Tc�sjqn�{%�*�7�*�x܎��? �qz��2C_`J�ݼS��[Q1;��g������G�pm���-�c����?z�Ə�k߿�P	�jG�Ѳ�����\E�2�>H��K����=�l��!1��a_�/P�f/�1�"H�FC�r0�����������9��E�؎'F�3��9�*�v�c|�=�S�F���x_p���ņY4�#g�3�3PD3fk��[6���]Ð)��U+ψ;�F)'���e��"����ެ���ms2�`�:�b�JI1�C
�+��	�	�o!d�e,n���������!����a8�oλ@;)A�j��2���9YHE��̡�0��D�?���$ZS�B-����6EA	7dh=p3��3�9��B)UT�Ps���yʭ���(,�j�Γɧ)���H��M[O[�e�KY����=e���[��p��+�֌ӁY���c�dsU������P����;-�Z*���ï�HC]�{xl��D}}:\�[�0,�h��#&�"χ��Yh{Zɒ�;�� y�|y�pnI��Å��ˤ�Ż�4��cʢL�uI@zM�9�_S�7w����z�M�ϰUGL��dx���P�!s�G@�X��D=d	�(�����R��{q�@%u�}�>���	Z�;İ�x.�H�����$X
ځ
����p.��(5t7�ޭ ��P/�⿳i�޵���L[/`7������Dw���*p���|� �5�5Bs�;S/��6��"x�;��:7�X&�����@�:�]4 G-�l��ĩ�g`q��P������5�dWA�7i����mD|�rǜ\��蝓'J����֧m�e�]	U�Օ��# E�'�C�O��e�������Q5�;2�������ǱV%�ɱ�8�E��93ȪK}���M��k�	&�P#>��L�(���;�-�ܮ��,�3s�BQ��.��5M��63�*o�'�JU�[]�i��#V��XO�����p����W�w>Y��Ww��՘6�#Tk5S�f�Ĝ�Wۡ3v�kԶ .��9Bb�=J51�a��ƝX�#`n\���o]�3��A��������tF-��2͝~T`��T�G�<�1��w>�)xx� _�4q��1EJC���G����'�]��ܹ9\Gr�DT��3Vf�5���1Bt�RWǖ�!\�ڰ��9�\~�P%p����)�&�\(���J	ȓz���F�_��u<�<`��/���uI�ؐ�,K��̵�Jς���̘�*�V�p��ޜ{n3�!����u�C�o����P��m>s72UM��Oy9�kˋ �M�?<�9�[+G��}�;��WvS��
!i>�1V�O�B����*�XS��I�$7���C�:�h츔h
���D����P�@Y/X��
��/zf�/p�ԑ/
�{����f)�X �jЂ�n���u��o��YR|de��9x�t.�l�R�� ǔ{�8�[-	=WT9B#�B�������k��m���b����iyp��B?�iܟx���tҋ��ȓ��)W���8ǒ�6b�J�}���x?v-��0�T�'�Y��G���*�6Ӈ�׮O)|H)�\%m��-�휹��b��*K����s��5��"�[6awcaO]�n���0�[X��\V�t����O���a�Dp�Es�ӭ��Ll�������;���1^ʄ�{C���8u@J�͚n�rGzͮ.�%d����ڃiF�K�z���q���v`�����e7T0V	�3�A�G���"t�y$6���)�������+��y<�+�}��_��ѣެ{{s�)�'������9��N�@�'��G��|��ka��
C�,d_S�=T'�S��n3p�6y!|oҫ�>��"M�	[Yx����2	�Q=��a*��q�(�x�_dG�ϻ�@'8�g�~���m��	0�n�8�PH�X_��RJ<K���Q�V$����=�.�MW��d<k�J��U���dVȿ�8�fqx���졯H�����F�kM�e6�̕I�F<���0����6uۊ�\o�*������~�`{E�0�D7�utm��e�o�Y�7��Y��/Nk���]g>`�*����߾�A�(E]��70ۈ��oߡˁ���hǔ��V�Y �1�˱O�߄���stH�أ3(53ETּ��K89���>���W�wɘ��"aǊ�sCR�DK;��ۙ�������� �P�H�H6MZ���籰tӁ3q^l�0Ԩ�m]] Q�-�q��F�|�oKc�����^<z �?\�+�T@;���TQ���W\���?���[/�bpPe��4�~=��+�*�?�9���m����&w�a�F@Y��>l(�3�Ȓs�'4�R$CC;�j�ҕ�6B�����Q-%��k��RّR�	��D;WC�҉���;fQ�R�ʼ
��,bh'5�}k5��Ϗ2����am'6��hLnR�)��i�b��Z �b&�Q��BH�x������D�k6��2��\7�u��Vm�zNI
�6�h�lj���n���@���]�%U�`�q������.V�'��V|��̝�A��$��O>��\�Lt=�����T(	W��Ptz��	�d��H �cJ��N$c�M�����Ks���$%爙�>��n�C$ﯵ�/�"l\y�"*Xn�*�&�a��2����8F=��\~L��scX.���G��S�2	�t����$�Țwٹ��
�e�oX\n4Qs���8PD���o�^����<t�Y֯�d���D�Z%`*8(LA�i���D1��E��ɧ��Z���F��a�N\n����E	AT�%�&�����(�ك������*I��UL�{�.(���ע1�&�-꫓�� �O�Q��؜ݚ��b�%�+��å^$g�U>w@a �F��7���������G��I�L�0�~{r����v����҄2�^�M<�>u�T.�x��:`�	���r&|��*�_^�aP'p�F��!A����6js�/	1����@{	�_����Tԝ�e�*C���Ԝ�v�b*[�'4o|O�G�(��(��Y��W�7SZ?����o-o���_�4�g�����'��!�m�O���	��Y`:>0��T���%A}8�1CZ��w%�&�\L~��-g��s�@
0��|S�b�0��`Y�ヮ��0%�5k��"~��,�sC+��s�&:���Ym<}�+�v���yY�i��Z����G3*�lMm���@���ܾ�W�'r�������ϭ�½H�6�q�?���/<ޘm$9F	݋��מ�M*��G.�F["�f��'b���^n���B��W���ˠj/���1��s�rp�ܻ��M�H懵�y�T��(��~�@o�Ϥ�%s�k��O	����E֘{ao�驦>�=���P4o�d�
���ޓ�փ��p�Ǔ�J�����}�#�U��؞+�d���C�Q�K�_�ҍ�A45�iΎr"���t���1-��5��I��ſ��g3���"��V��,�R�-�����	a�@�(�c��֭�4�;�l��J���O%����l����N�F��V;	���Ԥ}&"�M�����%������EM�yT���)���������U�v{����A:�!�^��!�h��<s�<��+����>�'�O�9��^?Z����ľY�^� ��9��DI���x㱆��v8;�XS���@#P	St��(���ucnl��0^�&ڧW�~h�V��	R���1j�A����|�qM���)/� �k�Rp1O}�l��j�����"��X���$H��[�9r�o��8y�W�Zn�@�$N���lV�w}ٱ�W}��Bt&��l$��m���2A|��d<�}GR(r�P?�� ��Z�����0}���(��W���.��(�_��B
s���X� L:�e�k���{�A�Qʶ�;��ĭ5�'l����(����j�\=���^�p3��qX䤿�$��'e�i搞�G8�I����e�r��U�'�P���F�n�D��2s��J��R�_�G1�_,��#��;�ɩ!�|�Y3p�GT�^�&��V���:	�*���Kf.;�׉y��zj�Q�4m��-��X�Q�<h��<��b��'����e���"{��A8Z��ugͿ��<I/�����U��\�:�܊�j�~���Ѱ[���q�*�"$d�r�e�2�qW�`�-&\�@k�Rҁ�a{��7W^�ivhv��k�/�O����Ѡ�1�PѾ�?�4Yzy�Pȓ�2WfXn��dN�O��TM*/��$xDZJT�"k����6:�I�� ˾n`Df��;L[Z�1�#�FH���As�`�+���j��f�KS���ŵ�z� bb�'�Ù�WpLq��ӇȚ��3)__�ﺗ_�����5�hkE�i��ި$��/V��vw�^�mB4!�.H����1�m�6r}���i�;dj�������;��O�z?ǭ� ��@�6 z��
Bc;T�}�h�q�5�,���y�����,� k%48�\q�}��żo�u����Ȁ&t{S�=�.y{��;%rKñ��{����.�:��]�z�H�^��	�֏9��s3�w#V����PΨ���RNz�'�+�ߧa�&��C
��v�as���ዎ/u%M��}�}L-�Ad�y|Ԕ��J⻺��bv�
1X��:�6��*GN��F>�Ǎ�j K�&�:��'�^dS꒕�>��Sڒ�5��/�:S~���L��!
�q�y���sJ'���+�6���r�(rI5C�U^	��c����5�X���J�^
�k�g� �rT>�8��
�����{�M�����oD=�eX;�w;0윇�o��or���\�Z��J�Q��.��Vw�#�UT��PT5$>N���Y�_�8��+72}�/��LU��w��A�OΜs��}�6�\�az�������[+��[�=�1��*�U�X���E�6��
�\K市�h��q�����z�>�m�a��ḛ̑�����}2q����������ɠ��
�7���Jp�B�H�;�?9�62T�nClﴛb��8����b���f�R}i�CsT;xG��y�~�+�7X]�H��7ny�*(_˭ׂ�钻-�������J��c�HY�:[�:�F���(ص�t����b.��T?��!�s)�YR�d����4�.�ﴦJ�f �R�.�r�\Ks&��7E���ϯ�Ą�5�<]���m�o������$��6���!RƮ:�w1Mj�z@�
��8(��~����"L��oO�z��V��������˚�Y�?Ɖ3�����9�6f�V��z.�Չ����ݭ�|�#��b� �f.�x1��>ʠY�3�errx#Gp[�[�0��������<R%�#�[oaI��9U��ۦ1NI�RR�O�Ψ�KSGG~��J��?�R���QT�ܗË�I����F�|� R���-�QeQ���"����k�L�5�fgjk��G��R������a�M�a����u�t�̍$�Y��a����Ϛ]��}�\h:�m�G�"�F'�0[� ���7@]EɈ�0��Aim
��n�n�Im-g�"��lX�Y�¯��F��)#y��\�h����;cHox#T�;�bc%�����3�n��Fʻ�i�x��[c�Yk�f��A"�w��Eܗ6�I1���~)TJ@W͊q�6��a~B	�*tRt����@2B��>�.��th:j���Y�������j�IZ�>A�MJ�Od[c��Q5�������0�H��`^��
���"�^�N�|)�˄�a{CD)-����(G{h�	~��z��r@ԣ"kf�1�f4���mԙ��?��I/���.|���3��tIFּ��
�ᰒ^������𫫚��9��+<
-�х�{����� $���LRR,������u�`�Ar��@����	��"=��2��9����
w�>9��G�sw�R�B�|�DZ� �5������+��H751�T���U��@���>�w~��"�X��K�a���>��+�	`ᯉ�f�;�ћ��a��)��.^%�˦@��g����"���:���%�ck�v��ʍ�y�<]��n��+
��ê�y��6��j^�񙷮���9��S�rz� ��v>i�!ag�>!>�s�����{�e��dX
�ʑ����.�r����ϝ�.Ŀ�jْab)��us?���G��6q��񕾥�>���k�ǘ�+{A2B>��L���oHc&��\��Q�U�Z��d�3���s�-�*Z�ƳӢ�|�@M�V z�y]���������zKRp�ȫ/�g쀁H'�,A���Z��~"Ax���q�أ}��s�k@�2*E���^���6��au5�8�1톰]p�O��2��"e3XOrn"�#	�d	w��1����K�Oma|�ޒ}L�V�p��V"!�c-f:�K�QI�\0��m.��C��Q��
JxiӄZ����n�㎧9u�X6@QP�TDvV[�R0l�'�p�I~y�j���M�s�ₐ�&f��%Sgir���C�H����:7��!S��,���	7U��=�o4ㅢA(Ŏ� d=�a2��}���2�>7u,h��%��t#u7����b'����p*��kʅ�R��Z�q���O��/4l{.���t��8!�4Y���}$LF��i�B7h�t���-'R�1U80�Qg_�B�!�
��)�#F���li�xo-����=����2_�*UR�"8v��F4~��Y�hO�:d��Q�Ʌ�nc����]~��N'WE_7U(7�'�-��cF�p�s��ea|^ȝɂ#~��P�K���3���o��kw��]�	���J,Wx_w5[Ż�����7�N�D�rH������_B^����%�I('j$g.���ؒXO2���H�i��ǟ�բ�9�8�����\��MV���������������Ќ�"p���\�2�w�tL�����v!�-[��XF��{YnJ��qr����}�'����f���㸆�B�'�n^
���5�[��W����Q��h�O���͖&��?��V平�8��u��ī�4�z����Ep&Iឆ2��e�(��<
6��g�Yh�������Y�Y�l��[2�ESiYP�� U�8fu����g�����D�o�����g2v������#���,�}5�Q>u�F7�Z�����َ���/�v㵥ؚ��a��p#7K����`�ƬwR�I�UInȠ�i��y�� z��z{SS��
�E,{9-�x�§���N��H�$���S�bF���鍽��<p|'ZGO���^j���@#�A�5Y�q:�h�A��@"���fM�$/�Nz���[��լ�{�$�ǢA�=̓�4n�D*L�]���.֓{�Ke��$+!Y4�i!�Y#������e CL��?;m�u�?t�<�6��f�+:Smq����q^t���v�Ёy'DF
�P�N.��-���)$��{��Et�;��UA���v�Pw?���YqYD�*Ա.�y�Y�,�i�\.04�c�Ǭ�F���O�s!��N�S�|;朾y��$�8<����9�x�@4����q�ܕz�@�0LX��8��!A>�҃�iA������;輡q�����>�K<�R�w��h�2�UH������������g+��y��l��&l9� b�W�R�B�TNr�S�%���+�24p��6���	>f=�W��B/]����f���'���>25�@�rt��~��?/>�M�t *����ߦ��q:�0�� ��msp sC��p3H��<x�E6�Nw���㺝�!IQ�
#����K�͘��u�rbX(�4�摱��J��c�JS:7��Bw.e�@&����[s�E3ϕ�KfZ8�:m�6C��[y+�z,G_��bJ�n#|8�@KG��g�`��2B.G� �I����9d�fL}8�x|scr�����植jX�=�+�ꑐ��Q&��RiH�
a�@��d��P0�
L�,�p�$���oqh��ȯ��/��JlL��w�������_G�$����ol��9@
�+��حe�����?Am8m��Aågѳ�@�����:��#F8nrf[dxOd��W<?�JH�s�C�9i��&��t��)�#�(��FfLn+�AQ3��jm��9& �V�s��A�WC}ژ�;����J�|��1���U�Oo�|��|M�R�I�>a���1%)�lt��Uz���*?�������&5�P��ycJ����p�2v��Jqû�0n�4��z(�o��`GDC��{f�x�����]�u�R�Ѳ��Rz�BZ��WJ�I�-K'�3s�Y�Bۨ�?��d������i"-�D#�Ԅi=R@-�c��������w��Ͽ��g��m�Y:��9B`��]�IR-6��GB������xa���c�)�}<"��[G�Ts	�v�Z���k�Zk��� ��������E	#(��W<V7�g�DMb�!��/ ���e/k%��#!XAxQ��U��OfZ���Ϝ9PEA��|;�;2��F���IЉ�R{�"���^X0�x�g��%���4u��[�y�xc�SE6tpAG��y��'�� ��x�BLv�$�h)@�[�C%zۻ!*��G퍜��X�*�����f�߯��T�E����,�_R�!O���$�a�s!�|�2�YI��I䬽��ڳ�GWl�'6��tZۯ�y��cר#'L�D��Y������ ����I�_Q!��@[h��@sYd���c�{!`ū�*��E ���t�&\���:�!
���/�K�M��Ԡ����9P\��\}yA��џW@�G�qr�+��ׄpl�X5K.����-���T��İ�ߔgv]</uoaL@���uy5�h���3�Z���c��e��˩ɳBzkwΘVz.N�-<���d��)T�.Ɩ\?Z�Q �����Q��4��e��_ia�[��5�c�U�q��*������s���(m'�a�6u狱Z��㘦o��K�P=�T����+͇r�uD��G�������}?Ɍ�&��A��g �<ϤL�h����������&Z8~����/�_}�����ɮA��'�(|�B��d�ރ�7�p�p8�9�#���}D�bl��S�-�K������]��̜M� �!���'��xH\4�s�3�)ߠö+�KLc6[ܾ@?jw �&�U���h�����~��k�<[�P(��Y=rr�A����0�2�s��o��}JLQШ+ʗT'n����ԡ�k�Q��RI�� 1f��d�}�����ο�GY��|��a���.������ƒ�Q��f�"A�ɥ��\5���WK�z���ҩ�9RO��0�.gX(�g�\э�(O��ȄC]t���� T�lZ�c�X�^��		��	�azh��ф����&���X���V�㌹�ܚI�t�]�nI3N驞���� yI괼���e�`rN�Y���w3���Q����'4
\:'=��}�qX��#T!Rl#5�0�xqVG�3�9yH�?گ^�&��"5����s���T��f��4�WG�ʇc��\��t��r=�y�� W�c�u��.CXA���qQ������%ړ�~�����`������q��ӝ�_kr�
u߾P-�؎�9���f[C�X/�6$m=��$4�A �x�Y�I/&Tqϐ��3CiiĶƮ{�jF0��o���O��fS�N��5W!%�	4�gW��E���(n{GY�rМ�������Ś�^%�Ć��
|�Jn�h7�|��xv�X�jG@���ŦC=�t�`'�ݾ�̫�M��#zȇ����d�Uv���h�V:���a�_���ٵX��L�o+E�G�4eWj����Lz
~�KҎa\Nb��s��(m�+j'}�y��V�[�}��_�p�$A��<q�Ă:M�j~����*���� �I9Mv|���i�6����_�e:��X"#F�n;N�E̔�s,�aS�ʙ��^,D���{�(����K�-�{.q���H>S�1�X��5���$��Q�g�pnkaHό��6�Vi�@�S����z�O{�SڻN�'�Ř1&��B(�R��G�,��P�P9Z��|�D�i����&�k�gг�%�����j���]s��ͼG��a1ǔ�`�������NVZ����Q��~�조�]��A���ӭ���)g�*�z3W�}�N|���ro�Jt	k�}e����iA�i,s�j�qCZ�� ��Q�R�+~�[��i%�1U̇\�����`�1����(�)W��;�( 
�3���p��9�؉�Pw (�k$�4����	SrFq�����J���Z.�=o¶�VW�oQ����Y�M} p?�IH!���/D��}ǯQC�V|W����ѯ�H�:����^ ��Y����à���˗/��L[�갢���C�G����٘�	����N{�	���k���z3 �/Z��؀��K��%D�Y����}�@Dpj��U:��e|T%�OI�,�9�9V_U6s(��I���͗�&^�,Q�Z}]���&����,�����zf�v[��m'<��h��s�?;���)i���9d���}>��| �R�����~����n��I1Gt*�O�@�d� �5	%�vs�6�w��d����MSC{����:b�j]&�����������g�p�K�Pp�XhA&��c��J��D̺�Gҗ�: �f�9��V#���tD��2�r~1@��px�H��5��o�<����>/g�����0��܃%X�ݔ��{�A�fֽr�X��L^�вa�U�X�KJ��d�j࣒�G]��M�%@�K$�
35T0�$T����OGH�}����J�)�w�gb�]v\)�C�Cc(�������d>���7��j��}ix�㱯B1�<�B��V�\D��t���x����%����&���[dx�Pj����S�)U��3�6ޒ���t��z[�D���{X�$�]�||���v UQ���%a��YW�3��_��r�B�"����Y4��ɀ��8��G�B�Q�i1BY��`�̉g��ϦBT�
�����'5�d�%�g0��_Z{�u6��B��ya����m�B�����A��������\�7�}٫d]2��J����	s�A�������SG�T�i�ӽKV�:!�	;�����ΑN���cLH���c�v�[_�:3b\ꍚ�s�k�k�Ç(��6��Bҕ~w�v6�����؟���L;����ntǞ�^ m=Ҋ����9IKLT�v�W��fڷw#���"�H�#)̐��4M���$�s��[i�����\��@wg�/�>�#�PUG�mN��K4��;Ѹܽ� &=�0�ϧ�%`�8�Ƶ����`����5����f�p� ��s�%^�|2o�B����� '$��q\���?R���y�&�(�'M� ���/�ϣ|O!ɧS˹,+��������1��Tt=q��J/���!Y�?�̄�^P���ϑ��:������5�m��*\�!�5 �S�[��`]���(��vT��;��Q���^�"����6���CVu�nҒt�����	�������V�B�Pݥ�MNZ7�zy7���P�L�My��x�L+�5��"n�%n��-��Ʊê5��mi\��{�_�xi�{Z��$�����{��=��t��DB�e��.��Mv�ԬIt�H�L7̞��	�����0n�������h�3���N�4ZmO!&-,��[k{5/�-�������(�Z�5>�e;��HqC?2�H � ��S��ihAzv� P[�'l�0��LT�3V�T�2���l��I�
�l��~3O:���0���/���N'ȅ�g���X�[_����T��Z����P;M�KQW��զ�M�b��������<��
E���wآ��=<:�rT���k�W��^��^0 �O"����i%k9$VyI�݆��w 6D����'�nu���3#J6~��yŕ�ek���F�
�rƀ��0�1���� {K5מ�=/�\M��S�p��/ZhNͭ��<�_�'?�Yi�+���@&Mc�+��ޭ~����"���
0{+������o���
���׳tM�R�����*�0 Y��v�9���YZ5B_������?(x�h��W_�S���!�[O3�9T2��1�GL��b��n�)d�T����c|��-)��R��⤵�φO���=� \�0Y|�d���x���,"� 9&�Y��5�ഘ�M�8���=���A��X-���V�w��bաY���qE��I���t �T)�w��K��b_Q"�IV'�*;�+���E�g+Zф�yo#c�7)60�U����$w����J�D=�,���>�׭h7j�&��q����k՞1L����%����� ���������*��	yY����stK��#�\��>��AH�Mwt�Te:~��9X��A�/~q^��v�8u�'�i�J����(�\$ f�AE����z��A�e���Y��ƽV��!������8J���[|�M+�?"T�Q�͑��4�3�8���h����uq�ʅ)]ڙxH���V�o[�p�	�����>|C�ʉ2��T�_�$7��|z�(]ɕp�tzq���1�1a=*�J�'�~����=I�e7·��Z~K�|��!$��D���i���[^6P�ȮtH��
�H����w)QIKܵV2�N��M���ך�J|&xk��j���9��txaC�x�C����CU�{t/S>��j�g� m�T�9��~�!��\�lU���6 ^82.�5׼W��U����ī	�
�s*D��"4�h05r0>X���Bc-n�)c�fW�>��
���p��]�[wgj<�
-����9Iv�@%��0?�mť���?��-�sI�$f��!�K�:�=���D����ls��`%$>�Q(�t���NV�2�Q^�
��2 ���G��)�8a����k��ݵ�� M=��p:K.8W���v� ��٭�+��w�%i�ˍ�����lm�?~�9�_E��Ryn�
>�3��/l����k�.��l�ɬ����t��gE�)���Ѵ�����T�v��^�>��/�&i�����:E�$n���GI��j��¶�y�܌]"�����v^	��'z������
ޣ<rʒ�@\���c!����S�w~\������u�:i��l,�f?����1�	�)�Z�t`��x�x����i��]s�U�t��WO���,�22�f&�/
K�qo8�y�X���O�̽��En���~�<U�f����YJO����!
g*�+S5WD>>��Ga�8.Hh#�5�����'����p���^��j3 ��1�Whs���$�im�{^`X2g'-z� �sTw-���J�r��* tf���������u!Pc_5ݪ��⫄��Hg�-c���o����BM�����3�T�ք��E��f���Pw�k���5*Ɨ$�NM0�ՂfA�@:*����][�P�Bf��%����R�m���0����ؒ�>4���2��$�qIk���@�`Lp���+�4*�;	o�30nq��$Kv�[
}�[���S�Wi�A}���Π1�O�)���i�� x.�Y)�Ԃ:��!'XI��=�s�E#��\���>�[Ήӵ���l�U�h;�[�Y�#n��	�=�f����),2���q�m�L��r���T�IǢ">°��8��ѝ�n��\�u���r�ސ�P䶮vq����^|�8�be\��(�����C]������u�|�0<M�dRl�㐄����,>��������MYn	�������|��Cl��MDZ�[b�Wl<O�u�'��K�3����ԍ�R�􆔥?H�X*ʦ*�	r�LNE��������=�$�%K��#X\=��c��*+�r(Q=��-���y�����q~m�6��ˎ����}_��5�&���~��A��%�/o��ʠ�O�~�/#5��7|[�\�ʺ2>����@�,�d#-%!���^@\��w�<2�L��UK���<�w@F��mYvµ���H��sg��	�b͓",?���M��w�y��E�GxEKM�89�;��)�_�K�E��G{�i'x�eF9֓sp�H������P��G�3Tn�ډ1E�z��2��vޛ["'N�Uf���=�`�Vȓ27���p̀O�x���N�Ou�������%�~��5f�#t=5�l����\t�r`+�rߚ�����Շ���F���p���7�o��م���Yny�m'��Pf���G��x|,��|0E7�#����;�\|ז>p#*P0��/ݗ��.��MyH%�K���ݸ
�8d�E:x�)4�E��e�n,0\�4�1h����rFe�z��o���#��ZE��$��f-�>�Wx�8����-0ߪz���Fd=Is:^����)\�O����vJ�FŲ�wɿ����t+������np��ڻeiwnh�s3�ÿ{$�#;,@�pi�Y�k�ݷD
���|NP���?| �7ة��1���,�Y�
�h�&ۊJ�9�j;����([9��։�����/��d,ƂH���� �1�ѿx˳��}�N��3Om��\����u�B��4r:�m��Xg�TR���v� ^Б6ҙ������������W&a������h��!3���XNZ����u�?��()R>�g8��	����b�!�vocGW�({��v��Uv���Ǹ�$��aZ%��N��*��P�2� 7�W�2�;y;�\�J�KĢ۶y
�lY��F{�oֈ�_�l\�	e�@9~���e���*��]���e�3e�M��&'��}��UPCA�oar`�|EX@ҟj�����<Hݏ�S�\���(�2J]�b�[ULH�cwH���Z���G���vĽ:r���D�Kuݭ]#5���
r0��h���0��J5b�[:D�>�?|�X���E�?UQ�T�� ��c���4Ёgѫ!㢎sW����F�z�XN��0�vm�+����,!������H9�[U������W�=��#�5ۼ�K_n�B������M<SaLҁ0_��-<-N�U�bu3!B�agq~,����8>�y���[I�mǷ!
>��۟L \�V���@�T�c��X���c�������{�EU`~YhЗ��5���; �FU �Kf�w�sŇ��C�U��q�u`�z��#�l9ֲ��,J��.���(s�bC�|̬Re�g�-�X]u�W[�ICl=Q��,��p#B��6�#VC��Ф�H��c5X�/g�!�#;���e��Q.dmb������3�u )+0��V?��h�1�)���;�iS�1</1�%4�yNъg���w�A�JC�z�6�{}}���ǻ����-g�}1板0?Lek��J���AVD��Ԩ���%tdw�X��2� 6�\4�|a H�ȃ�f�݆�,Zܞ�u�S\)��/}a��
�c���jʌaP��;ڝ5�s�t�����g~�%F�6��@pӺ��O����7���x��C=4�	��$m�)��B�xVK�y����\�ǉ��7;��*�?�V07��_/�ȓ�C���`$y�_(᳝�ÁT&�u�	�q��h̡d�&���}i>>c�M��f�ȴ�P�ra7Kk 푕")6A�罈��c�������63���.=ܭ�f�������;��.:R��w���6B���VI��b�l��7��.�v�X�.	�����XUס� T ͣ�gb$:�����.8���m�^�{�Z�ÙB���d��U�����=nH>�{�[n����&_Br�L���X��C��V��I�3�-�BF�6?I�?0�/�7#A7|)�Yq�Qe��#�Fn���o(hZ�O�;�Ə�2P��C�."�R��������]�G��4�&`�c���z�r[�@����MrP�1�.�@4��h�W:���.�
HkR��>��Uȃ<vh���
�%�R����
���s�sSwb's2��X#���*=ދ�B�m�E�`>�6�/OG��2`R�Iʗ��ot5�8T�l7Qtf�˖<��O(�ԣ�{�{ͭ����8}g�\0rפ��
�|�>�C�.�¶��e���H���2F�j�#9�6��n
.���2����Y��-��
aC�u�BПk�|�](_Q���Ǳ�U��#�r��IM��p��w�#��9�������M��3��}]lځƆ�����75��}dE��(k$�ws��B�i��٦S҃��lNW��|��>����6E�>��ఞ�>P�  ��ʷс뭊�A�8���M��\�Z�(^L�hbC &��S9����ɶ]h ����7{�F��<e���Ǉ�4T��lJ=;��AΨ�t��@4��e�W����ڑ.f5�A��Ƥ48]}�}�H�����ɟ�$r����6ZOZ"JM^�*��ՋOw��e�0�:ZGÃ&5@����R�	 �'���l�d?`�O��V]
����~����B�������ev#�iSQ֓�6��Ja�Lm��`M7�h���;f<6u{��kM�;�<�J�Ϡ"��%,��؞��l�.��r�i���X�� S��W�B��;��K���iM�-�#�E�i��L/�L���uC�$��̿�
�i�IBw�&85��1�kxk�(�0�M�\�B��W^�져&P���qj�f�Z�.^�yp�>쉬��m�FթUveE��� SȂ�f#�2>����"�&�bzb����g���Nfd���k���A�^��4���K��Ga�;�G��Ec�g�70q����E�f��;1ö��F�#�fw	��<���k����:C�?�ňw8�X��k[�ߕs��wo7b��$n�a9M�F�]���ˈ�t�ֱ⦙���Ϲ񩃪H�\�p���,�\�'�P4�4����(V�+��k=�\�կ���:�׃�T^����c~2Js*���X� �3�&S\����Fd�O�����[���|`'GJ�c
���j2#���N܁���U�h9&���y��q�-v'ZY-�0+�{�b8�ߕ;�`����j=Ș]��r��'�sy#D�Bma����xT��.�>tRΰ�t{0�o��
�($�Ru��m/�m�ՂNP�
��`�o�EX hHr
�t|n��
��jYo�<��h|��۞���=%���5wH����M/J�(�84"�M Sr?1N!�"����O��p1�Ĳ��r�i�!����&��`��\��V֎�Q؎K"�����3 줷��T�G8#�3��;��`�"�_�!"��؏%R{��X�}�w�Y��)zM/	��sTj4�Y6L�� �,��2�W�H��
(�1 ���aN`K������QQ�
E���m�D8��r���܂�����+'���-֝���_l��ι���ێ���WC��[���7������`�X�ܬ��k7[�?ȰHy�����n����#�ĺ�'A̞G��r��N��M��1���&��S$3�f����=���õ���:(�8-\ȩ֩��L�d'���vKdL�S���=!���,�u��!��9ȷ	5�ͅ��ⷔc���jY���?�jצ���Gb?���s7^G��}UXahN���,�� X+���S�_���=	kb�/}d���.YF���U�]Ls�z"�>�J�q��1��- __���Z"�t�EL���I����p�,�tkY���J�$�i~9K��ɬs;"�2|����Pnn��łܟ���Nϓ� K�_>�s�T�䡈X�{��w��'Fm���ΰ���I}#{�J�b�1�^��V����h�zw]�٩8n��$�EЖV~��2�6~
�_WN<%�'Č�����b���Wۦ�#�c7UBW�g�IAE�#� B��goA���0*�p�^]g��9h��f����@ao��E��2O9`tf����N��Pb�Z@�	��'��j����Ì<�t$��K�~�����er�Jm>�[���c��6c#T�z�q�珩�C*��Ƹ+όd��D�������«2��3Y� @��4g���DvVY��R9}�Բ�"�0<>B�9�(������6$�f� w7ʒ�Mpv�w����xЏ#�d�� 9Z�<o�Y���&�I���~����>�gٓ�SK��2.���,����?�eVMO�>%�_����L���E��z��#ґ���̈́�`y4#��yZ�A?U�O�fƒ�f���|��u`"V��z��tX�Q��Ǔ�k5���^5�
E����� 6����-v�:��)��C�S�~�gæ)A�p�cԍ?4yd��"�4PY���`M!ns��WzA�Z�w� ��~�NWGL(�3,�(��ӵ只a�^�;�'h��l��EP���r�F:4�c�߬q��,��`ϟ���z�@X��*��+7Kd��o�|� s��1�-�~*�I@?���[�t�1���1�s�D����N{K����r�|FCP�4S�^q�#��1#����Ԕ�@G�
G%	�6��#qkn<i������T��g�R~��u��76�Q*�8-�!ҟ�J�_�&�LB��`k<�ۧ��M�6cqG�ѩ�7a�>s���V�ʌ�?�w Q�W��؟���U��|єW�[(B�߈��e��lu-Kz�q������|�^�2��^-��몄�p�D�RCV]ӧ�O|L`-0��g��4��.��_��6� ]zS'˂��qnM�p��ˀ����I�w�K:R�eg�sy3��a�A��(�%c՜M��+k?,��.զ����7���ˇ��C�j��
��'�6����C7=:��}��0�?F��+�u�W_��II0k0}²w�)����j2�o���
���S�٨O�Q)uJG��Rs ����QK�e�ҷ\��߭;�����TL��ȉ6o�-o�?�G|��p�f&f���T�;�C\���.0XTR��WFH�Ѥ�֕Wo	J��j(J���?一;��6
�T+�P�p��Q��B7U�%��ޗ�m�Z���Fܙ+��o} T�"kj1j��a�{�H��k6@��;���	�u4���n�"Gb�Ѡ� -1땼�p$L�l��ᵅK�QF��AY�Bm
��K�p�V�2D���XΡ=��`'������@�iI�}̸}��ZDS���I�W=x�L�[�jyH�tb�#.�mA���B��.c�]貫�_S�̫�d^{�W��{"��f���f��}�yoVU�8�WK��������ي[�?�,�����s��#-%r	��c���z4�ܥ��}Cak~��H|�7^Ff��GU07 (� 2��[��͓��~�#��H����BVx�3�5��X��+A�ޱ��!~��hH���p �n�]Y@`�f�t�'�_&<���[g-^� �LA��̗�z7ܐ�|�e��ޥDN[maMg���ݾO����Pv��P�w[1�F>h�*�#�t��p4i�/}��I�++����bCV��,�w��y�q���R�3���ƫ���n��,T��b<U�(8
��tᭊ̑�25Iw��wA���X�y'�<��r�Cw�g�ЃֈC'O�&_ߛ�r����X���}Ѧ��p�y/��]�V�l���M32?~����ޓ���Q��먃������'艙6����ՙ�9�$�n+I��)-9gI{6hL"���<5q̍}u���F�7����xY顔���yml��q��#��a+��`+��QW�ʾ)4zV�Cq�ԕ�e8�	�H����Z\t���R����F3�p��a�t��N�5�Iߍ��E���L���Xs2��@ɮ����پW,#ǋ���Ơ�zn*�x���?s�8�u+q�2�@�H6��5��2L������l�FF�P���6���e��4f��sS�-���q��7�C�5�=,�S��x�������`�H,�$��yQ%G��ͬ����ڻ�`D�-�g4m(: 
Z'|�:���V.j̞!v�Ό�3�W�q!!���F,�CD�1�bmu5{dJ�,�<��*y�`�P�mm�
���韴�rR���YG`��m4{��p L�t [��N�n�v0��D� qۑ�eb�*G�I����C�,QM�y�|_v���,�_�f��c4��҅����j��	�- ���J�;�^pM��͛��FX�ycv���j#PP�#G<�z+d��M��88E�}"+*骑�>Vb^�K����RP��h歵=�fa����{�݋8����\:��|�B�L�n93L�8�F!����~J��������}g&r��18el1��G���-��]A���BF�N�p�X4�����J@�|2É��Z�ը 	��-`��_��kj\�HA`R5�A.��_RSP����o�����`V��f\���o�
"�p/1�_����Q��E����ئ�u�>
Ƹ�!�9ǰ�@$��u�ENY�WMRZ�:�qٰ,��5��k��
hn�kq���\:9����ފ7V���b.ɴf4�s/������Hʑt�zB�i,MO���@߁z�h��ؙky$��t	^棁3� �A��Ķ��z��b�>�c�T��x��o8������|�={�=D �L��H��~��a?�PqO����7w��icd����ru%We{�Fz��RS#7�$-���e�
�b}����p��m�=�)�
/�V��y�m$�8n���LY�Ah���]�� ����[w�ס'��$H�A�	X��}*�r�5�X�mĊ��G�-��������&�� ��|��i����{��-&:�s &���QН�b�>8�o�+ }�:_ܜ8'�R='���'Qn�?�E�>	ȗgϥ
-Y��j�2��4]Z�~�&�R0�ס�wr󶫡ng�R}�=���2�&�c��L$ �\q�j,_n򅀼�����(����F��Hb��-�A�ʦV��Uj���H����&Z�ϴRʋ�p^Ҕn��T��9�KJR{ rϐ2����k�`7+X�y68��ad�"�3�\�K|�2�M�������eY��i��=�y���V+:C	��yr�suLyA,2��H����o_R�����Q��d�0��Z#�����9��J2Gnz`��K0���j�_�Qs��JT&{��b+���ㅏ 
L�h�Uhy Q�ut�|D�T$h}_"�Q��5yC���d���78�����41�Ͱ���uӳ�&�&����^?���HoN��Y9�V�����F�rr�_N��s�0_5�k�JC��݁H[_��r
�⦗�k�0�꾊2&Pp�SwRɵ�t��ǡ���dMH��w�͟~���;��ݕY�Hb{B�1����o���AL���.����4��(�6
/��_�K���tɊaI���y�^w|���Y��w��o@f�i_6ś�~�!�����{
����ف�=���}6�h]aF߿�$��Y�Nq<��~w�����?��{oe����A0�d�u��ItL�'��\�S1����w���,��mc�,�;U`a��T��JKĴ����s�9��dj�u�Kt�����<�{��+ښ�"O�����7k��P���,��1��":��O_aDo@�ϜU�k�Y&�|R6!�܈���;���E�;���q��O��:>
@d�c�{6n�8�`9��̆VK��;����9$'��$ܷ&�Q�]��(R�b�S@u��k/��'*�7����ߐ>I^�+���Hxm�����2��@�Cӹ����I��u�%��l�q8��r������zō57]u �qߌ�����Z�!�9���P��l���G�L3�w;�g�xl��ʈ�>G��'_��j[�t��D�W�B3��:�h��"���hq3�&�|�\�QB)2��䓿�2�1X�w�2~��D�����^���̮r.a�x�-��Z	K�v0c�Ы�u�O�dƠ��B��#�)����nS������������ D6ѝ�U���i,� �X@�.<�
z�ݕ��EB�y��;�p*.m�|���NY�9��b��3׀�cdˀx�H�r��$p�8_ �+�4�HIF��{b�������c���Tg���������z�0
#������cL����,O�(��
E�`U�+m�i��i�YZH ���zC�Kv��F��n	#���-l��+ɨ>d7�1�R�N�)�C`
}�w�ɝ!��`2a��T�o3��b�G��EaDJ-�B����kbR�jHJ�|����N�L:�g���%�BwW<��-;����鱈P7�m�K=d4�v��]�5����O���8��4�[��f��ȓn���������+{IXB7M�Ҏ�<7�߶�ֆ3lT�����?��D�f]+���K'���'����vs�?7�D���ibu�lַ��Q�я��>�E����(�<��TvN����ҟ�K��ep;���"�A}Mg���V�edjb(����� �� #`(E��Ju����3�C�G�=X��A��>�ߑ��S˽����_k9N��
��k�f�qg9y�N��s�t�ō�]c8�mG���"�#BU��n�yd�/�U���@��Z��,�fw���6����?�����/�����񝖔nz�پB