��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�?u G���F��FN�t�����<y�l9uK�P���+���ú��Ŭ�5[��[޹�����@Y�]1͏Y%�7]uGq��h�ʀ`7��N�O���/�_�͗�oyd��4�&F��\���`{f�j��yH2_�C���b�p���'S��Rv��6M���ǧU�D��r:c��Y�`c����8y3�K"D��p��̯Ն�b��/��;��]mN̙�m��`S"wb܂��l�@-�x+c�v�A}����U(Ꮟ.2�C���Sg 
���8��&"�<s(��=��ڈ�t1�ګ-���7����d�W!���O�F��<D;Dn%(ZM�&O5�*�0�Y���]�v9���.2!���؛��.F����h�,T��yC�L	Lɇ�w�+�Ws$��rs�W��"%�4���#������J�F|�)h��{����Va��j%�ǐr#)��Z����W���Q�HvP�O�Wێ��m��Z��P�r���eC�{���1pw˰W7�X|��o����o<�
�./-�Y����ц����[�Θ���h-M�꒭�䘤Pbˠ]0�N�~V<���ފ���5�Ht�\(e�}���5���������Te�9>}�p� �"��Op�!)_ ք�d�y�D���47&70���x�|�H���`Cl p�����SkD[M"�D�xk*�!-�q����X�G�|?�.7�it�F���G<�2��WHϐ�jG�����,�#al�$�bڀ�� �L�jBΡI�!��Sd=N׺�L�v���f2�0I�8���ԃF`Gd�W�c�+`��*Yu��-�j�l���/;F׸Y�=t���̋	�)�~�L���0�)�0?�,G-�݁��㎦��H��ٍ�̜2��tH���Z�ml�,u�I��my�`�����z�̓��ń���*��	z;�]}��j�W\A�csֺ�Uμ��F/�?�|��9��������Z0f���y"lq��@E�҄�+!	�����	��U���K��v�y��N���*TEt��Y�����U@~b �)���
���n��JNg��[���_ūt��S��r8�5�2b;�z<_���L*���^��Fܽ����0@�?`��{g�����P8�Y�Qw�{��O��JD��b!���-=1����P�!:L��S�o�j� vVzi�y�Yb�d�D"�S�ck$穒lRO�I�/��|������g^����0ΤG	��z�M(Y<��>��h#=��a�}.�����u����,��~��(��jT��?7nf�H��5ݭ�0��j�1C��<�#}s9�����>ʝR���P)��%���cqE_�s�o��[<�5� AGfp��}��wA+����P�[8F37bB�FX�2�P;6�7�[�^�v�~DUc��>��!f�pZ����� ��J��7u�2�QbJ��ʟ�]��u�������e�蒙fu��ͫ9�����g���lM��DfmxG@p[.�����OEҳ0C���W2�u|`} �gRݷ���*9$P�HFC����Yi�"vϙ�VpPk��ђp�_70������c�c��b���l�5�O��:.�^	�Y�GB�k�e�}A��(�tWC�1Z���T��>�˻Q+ 0��_���9�!gB�D���9���`V�����]��*�T슮�l��l Xp��3�J\���CA��2���k�W2��:d]峆8/�v+Zؾ�T��� T}�7]��'��J֢�϶�����x�'*���
V������M"o�֣.��H��F��8��,�[衲G`߉~�$:6�p1���
u