��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��v�N�쪈��%���ieLF���z����$O�� �I?�r胬���TeUͷ���ϴ�I�'O(�y��jEr����د��6�P��y���1K�\�4ۜ�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�i�8����!ׇ��,�.bv��.�$��-��ig��&���xg�� �ea�p������MA�E@��ӬL�r��z�k�6E�5^Eu��#	�W�ڕ=�v_��Z�H�� ƿ���^5�Rx�s�n����?�R�����5��D�V|t���y]�q�Θ��-!߁_�W�.c�!����C���0�z�i�H��֚9��R�*��� �A�Y��>{X���-�^�/����*������P��5���a��������NwK�j�k,(�����. /�8���	��̾�sx鳽�=����Jct��o�r�~�>AM���
����ы���-�3Ȍ�4ſoS�լ�z���%��1l�18s=�$M�'�������m�����U,���b�4+N���u��T���n߫���VYK�6h��7�Ջp	��^i�a�	�E� '`�������>ZH*U8mй	��^a��6�-/�r�������F�c*�h5U�Adi�>{��Q"柦�i����Wk4zR@� ���fWR�+:7!�B��8ωL]��\�r�@_CE�'(���i�r0<.����\���1O����/���	p@�5�����-ۤ��UK��@t�����-�s����z(�7��Ȑ;�?�)�w;_:�>ԁ��A!���D���:���w21M^���F�Bq��(�� z��&hGS���i)p�A���+z�Rbݮ�sû�D�fd�.!�C���F�+mb�.�-�3e=��U`���D#�|)�he�����i�E��*�ʹ����4^̔B���/������HQ��ح�㞌O��/[�D�Lu��ǲ��Q��A9������rE��|�:�[�j�o�	D��{S��n��>��кVgU���HsF���l.%�E!G�d��>Î���h����7�v͠:�*�O��V���� �{Ġb��K^�#+Sh���,ǋ�咸�[����8�؁?����N��|��}R�U� �`�$�(����bv��B����m�[#�lC���e��j:p�y5Z#��86�}�)� ���X6�~�O��ow�	'΄�9��x~AVy��[�غ7�0��o�^�O��Z�{@�Nʃ��\�uY/۷'���p�}&r���:	j�^tN_�����fl�fk���c]~;���e��}��]�2��"f*�6�s���i�W�yއ{r�y$��RT6���35N����ljQ`v=��&���1Qл����\����_�?e��l�ȷ䇱jz����(��l��˄�c�(yfէ�����/=I�8��hru�%���.����ŏ
.��ֽ8=�#em��T���#��vT@~o��<�e��qϙ"��d-����"�+FE�ϋh/_�:��"nW��9G ����u���e�H2�vUO̮�v�?O���3X��BL�����xz����xO�륷��۱O���w��Z:>�j�IBJ��K�s3Ө/��{<S�͗�9*[������ ��T��ȣ��cc��x�J�ȕ$���E�l��<<�B�֩�c�d�b��,7V�k�u��8]1����	����j=�G�����'��$ѭ��U��
(�\�xȩ��2��z�u}�O��+������pck�
�����k��ѣ�dz_OS����$hQ�p0�*�kvħ*�0ƥ*G��,2����Bi�c���s�l��^���^��
�>����MyK��>)M?�ҴR�,g���B�;�d*���v�����6-Ja���͆PF���+A�9s�f��9��_���&>F�Ra�	h�0�R4,�JQ&�b�{/�E$�W���MR��2���x]:��܃�f_*G�;�?j�r�a���2+��yԞ,$!�(�Ow��aH:����x�fy�^����%��¥5����E���|��9uh���)S�U%š�F�{�\���$�-�.z��[�k�yTE���o�r�u!�����"q.Cv��b���A��s�H>�j�{�b �.~j����8AL[�������g��A���b��S_����3@Di��o�����!M۹�E���f
��"m�]%R�L3<� ���u�>�z��j-�I�km��:�UW�xKN�~�7�'K�2���iYR���k�H�����ur���#��!��P-
����0?�S�����L,_��Q���Vv��������1Ք�)\��h*��@{~����(i�����^��]�S���➯JY�䭱��Z%�����0��m<��q��0i��o��hf�PNv��S����gf�*�[����+�t�=k�-tc�=��0��.vF�_$��
ԡ/=��{�lV�p�!�+@��<Г����B��}���k��x� cw�k�L�����^a0wL;�*!�K��,)F6��� ���FI�F��:6R�
�Yp�'74ܡuX��V��g_�)�^�)��Fe���dh u�|SB5w��:���b���`����v0���ԼTsa3���R�%Q�n�m�v�c����p
��X������E�Gt��dK��,����i��҇�����$�y��X|��J�Eu���P|�>����\ˀmLϨV��Y[$�~L=�O֟3��!�k=:�R�!V�gdmH)��)Y�@�v�-k�k'$�z�=�<��2��$
@f��i1D82��q홒H�e�!9<�P�(q�[�DM���T>�ͣ�I�{���3�H��5Э�Gx}�-���vR��<++𨶛�"V�Q��Y�)���a�s}9��:���=��Fd\�	&�3�T%;#9����y�]�y)z�s�K��0�+��ݝɺˏ"G�����BІ������k+�>�P�l�ϸ,EQ~�ED:�i9��-?����C^��r<����6:�/hwZ��Z�2�2H`�mL�����S��K�,6Jԭ�%�����9�	�ө�.��}V�&Xkpv$��Z`��I"����oക��P�>�X��ܡ �1�g鐮�oh��zX+P�[�욾�^�F�r�����!�zX�0�M��|�T�5E��3���^�azD�ԏ"�����4ݙ�)�PUkx�ia�����;�|��{��.��@?��<M�JwAګ�ρin���Pz�,.���Z��h��!w�r+Ġ�G4�� �ƇJ]m���Wuh�����B��%��_fTM�d����'zx��[��$޵�����A�1����F�m0*l4y���8���U��i<y��@�v��b���?Vv�a��_��Z��-i	�����@�v,��Y��WA4�5_���u ���kB������ �������Ӥ:t��^Z�Z契V�bx_�((�5�D������ʦ�T˱Gu.�?��P&ŧEGB 7ހ�{�đ@~��f5�L�D�&D�8H�)�\}���DK[5�m6|X��n^E-�(~[E���m���,�H�6�[��&!~�O�1�O*���h��֙Yg@[I��w �5Q����0,O��Ws"f9y�#?���OK�>W^(�kC&�I0D��n�q!��#�\s����a��{+� ��+�J)���D�c|�p���⮊��N��9�C�޹~},�8�7}o�DY�~=D6I��L��S�x�] ��=�e�V\�,��p�<�Z��h1
>�Г�G͜�w�ό�hɊ2��t�\V���h���y�E�/�"(�Y�f�"�ӭDy��¿k_�y�z�?���o�\?�g��e�L�4Ú��Բ"� ��h��]��z˽�����j�#��1D��oN�#)�M8�E]�@����E�����_���p���1�Z~���L8�I"<�>s��?J4:u`���?LH���'8�΋���CeRkL��!��J�8T��ۊ�n�,=~q����M�h\p�v*ҙ��<�v뮧�}i0	� v���iMk�*�9t��!��b�=
�D�����&�C��R����`V�4��p����إ����ATc"t�t�7�<�w�ʒ/qٓ;�{��ȾR����r����lZo�p:b��![{�'�Q��ҋ6 ��h��lu	]��k���W<5V�)NZ�]lP��1L����1�HՍ`�'4��r�Kk�B����76���q��;�>���5�&=9��fҹ�i��6�>}q����(Z�}Ln�)��#G��˜L1��{'w���ʯ/Z�Cy�=\�����.
���1��ՙH�GA)��L��e��u�G[ Rm�Gc{&ڎj����a���q�U�,�a����*��b�˫���l�'xU�a�t5��Ǉ�����mY�R��ǉ�cYEӢ{�����6�8�z�0��W�S�)�z+�U����a&��X���ޓ�����MDJF���kTs�n�4�%:E0��Zq�����{�Wf�$ik� /0ͮD˥X��0� [�ōl~[��;�z����Lժ��\Y*҃t�����\J���Y�{?��fz8Mϑ.e�[����lr�D�5DS�y!�g����c�͇�j�l��gp�Q�A��+3b�
1�,�,�S�iϏ蒌����3S�r-o��\N)���ʫp �.��-�p�o�f��\!�х�������rY�F{���F*�8xf7b��?�	�y�vw��Ѓ��Mړ�m���v0�3�k�Y��
�T����P��T=�ˆ��3�ݱ���&�d�� }aYȻ�;!L,�SL6�� S}i��]5N���$�����U�0G�Į�5�1� �\U2��D�mc����wHRɰ�  ���gb�n1�=�3��rEu5��W="�%T��m�W�#�w��N]쓋ۤ<�f0��|/������J��
Vd�D��'�8]�����'�f�����3-9����+��Q�=g_��b�R���u����DVܥ�AS�аFݞZ��_9�=�p����j��V���^��g�3@��'�(��7�!?ܨVg�������id �fhr��c���$6k���JQ��_�����{�Ĺ��%[z#�o~�_�L����(9��^����0�/��#����`�3~`ӔC���`T 
WI�W��na�df��� /���;3+�e�M��f���[��%��&E�:5��#�9]+�u�K\� �A���荝K��ge	k�K�'Ą6ܦn8[!�37���cd�*7d�����]��^H�V�L��7��cʅ�<�y���d��2_�e�����Xǝť�
!�R��qg#Se��~� �?Lz޹��)9�	�!�����:�w�2H��y i,?<�=�mN��<�3��f�
�Y!�d���T���u�ЍS�AR����8�:���䯒�ɩ e+u�&���}��)q7�-w�JJ¬�����fr�"+�1r�;�$�d�H�9�R���� q�����F�,H�p��+�ж^gj,�x4����ܧ���� @5�[GL�ic�+�����@�����
VMN��H��C�� ^)��c��hWVE0�A^X�b�"�q��Ca��9.Ǐ��jٻ�1}�H�՜�sw�mv�0l�6�8�N/hGώ���6���Qɥ�zS�,��L:���Y7.+z���˶�3�4[}Ǽ�N8�'2���_a>�ޜ=G��^�8��rc� �HD��9/y|ɮ�qA#�����+�咅+l��qH$�|>�E�U'89.?�&����^��c��q��|��'4I�"Ms�*�����n�2��Eb҅�[f�˼��W�h�\�_/��`��_�a}[_)V�9��'��&��1{g�äd����c��j��>3�]űmڝ�,ߕc)W���������1޾�}m�$.2!Y4��?�D��Ne�|I�(�!%���v95!�u\ɀ7�PLD�%�c�j�[��_x��#�N���i��l	��{����N
WW��5���w���6�V�~?`$Ɨ��7l^?[JHUt0+]�N��Ф6M6���N
��A���[����x�\3u������R�w�1�m��᭄=�&���rS�:�%���قW��@.J�爫3����{�&���Eا������[�>�f
��S���Ȝ��^+�}�q�L�z=G�s��$9�T��j
_7	w9s�LW��av�ʏ0-�3x�眵X��oze'��/�v+�V����H�lgˋz���Br�$�$����������$^c���.��e��[�_�~� `�bK_jSx�5��:+�G���&W7�5l_}��:�M�.ة�4�-Q8��浐���?���%M�V E�@uy�H4V���PQ��������g��0��nW+&��/�2��ɳ��-�͸ �NU�y"�!P^$���>��R��o'�9���b$��F��M��Z���u��Z e:�&��w�Vp��a�qa�=U���W�CRZ,/-��[�+�D�K�_L�x��0����I`"J��*`��Qf��j��:��(N!V�UOy��ʤ7T��	2l�*��R����O��XQ������)��wV�Ԏ�.�Q4j�.[KXzb(39��E|�{�7�l�!f!e����D��)�U�"�uqY�{����ŗۉ\4ٗ�1����� $��)��ٰ%JA��l_:0Z\��.g3B��Õ���1�=�c��cC",,��v���A	��bs�J C�;�Sv�G�(i���Y�BX�;.�B�˩j�O�3�����#([3��6�+�+e.���e:	Ʌ9va����7���Y&�a�*�6���
��m�����8�8<΀�/�;D'�-��Δ߇�>�	���%K�<n5�)��uKU���kωf .��\n�Sz	�$r����q���PP���6�+P� �������m��Z��:����T}אټat�.Z�w���orU;tbO�}��*i����8���V��&ە��̹�Ʈjrj��mK�Z:�����=F�H�m�| ��#FF�G��M��m,��dSǐ�@8{b:ڱ���ó�Ĵ��w�\;��l�5��2��+n\2a�!s,icyn �2YP�3�Ϻ�!��aǐ��7���jP*8��� ף�@��d��r@�0�]����y嬎t�2��\n|��|+�Q��_��$�^r��Ɍ} �3��#Z��K-+��mM*^-
����K�x��?#pZ�`�!��²|�I��R+V݌��>���ni����bvNJ���$�s��)��{�Ns���ۅkn�3�#Qfr�C7����8i�\Z��Ƴ�����T�U�[9r�/���Qn��~HrN��%��F߶](O>���&���Y�!0�c��I�Y�:���i�M=`���+��!;�~P[��*Y�a���O���է�XY\t�+�;�1��,,:�������� sED�P������y�/�w_��䨫zH^���r���Wp��U�{�K�[��c/D�j3��У_˟������j�w��������|bzi}���o��7��v* �Xa���:�y0��7����LF
u���4w����=y�
�X��OԴޙ���eP���g�g��2n���{Gv}`�=���A~�`f�W�����[�7:�8�O��Eqk>������>[M!)X��w�똀Ē�d�NA ���_�j�'C|��c�q�pX���l�v�Q7�w零W/�rd��[Y���@R)�Z�ͭڹ��Σݜ&�`�hYA�׷M{�O�^�+�3P&�0i!�rԢ��4:b�L�f0�8q{�"���13KE�'�CO��[�H��^�$��u$Q-g��^��Yq�&��)=��ys�V�#g���8E2��%q3������Vru�6�&?�"D�č�JiM�S!>�=@ <�����+��b�/!���2�i�i0m�لZ��N�u��X��I�M����G���]b`�H�M����n֙E�a�|=�c��`��0����No�pZ�^���NQ.K��X��{N ��%��s�78d���[U�L
�	M<ml�x��x��'g����+�բ����;��t����3�o�{���i��i�,�[Cj���yacJ�	Z'V�M�!�&(ը�����D<4�\2��Ѡ:�"�`�y�O�ݒ�vY5��/��`I�R;̬���?�EƂs�쟟(�>����ﰚ1�J�\��
�z�{Y9���>\+~�����V��{(b>�fB�B�[!^� m�``��W����8�t�F�����DD��f�U�鎟�*��� ����w��-=���F]��	�"b�BĠ�%S� ��ؤ�~��p�����:�DI�&�&�0���ɕY)O�fb�(a�ꭠ[�}.ה�N�HP�	=�Q�J��
&�V��x/_"0���)8�YgpܛjZЊ޳ o����ax�Ϊi3�e��ɑs;b	�SƧ(���3���c�������=x���v�
4B�Q��I��m���b���H%9����ŏ`0�W|�%%�&4b�AɆ"��4�I�C�*[�`��습`�$��'�b�b�w�(`�a�Y����ܚ�\�����B�ɼ�;�uVe9�[���1��:��GA�R���(,��;8��Z	�~��˴�۩qf?��Jq]�xys�g_={���ǥs���6k<��/�om�!�eEG�iT��-r-�	�?H�o&���T �l�N{����������r�oA�	��D��ܕ�� b���x�^L����E�Χ�9$M�_I7/p"$,'�/�v���4�Jo��{��lo�>HYZr?�/3�����������I=�Ctò��zp�0�Z�d?��^O�0�����Tj=�������1m���ܭ|9h_SPv����黪=�B��q8!�i��=� SI�B7}\�����E��hR��BJж}��	��&YKP">��q�$�k#$ܒܟa�U����?�T+HD?+�2�u��Kb�-�Nh�s���:��η�M�W��$����(x[�g��Ϝ�G���q�	U��m�}$s&��x"I��l>��ڌ�"���: �s+AgH����xw
y��*2���z�̿ŝ��JL���5���>- ��]s��X�7���f�jF�v�uR��ɧ�"�n�c)e-�?A�3��S��c�0��.l�i�7��3g�1i?l��+`��|Ι.�w�F�pTy�fu"���KF�'�^��љ���Й�`#_P1��V�K��xL����"��W8/ ��Q��";^��ޖ\S�^@"��i��)?O������	����������l�F�x�SSu#�Bר{r&��rzZk+���@7�?[�U��pH�6I�Z�%P��0}	����j�ט�Z�Y;@n�����'@d������l��*G��õC�&~�7�ȫ���=��gD�U^�%��T��1J�V��!�9�������o{!�=I�$P�'$����R�q��f�	[[3�M��<:4�!{�+6Q�,�>iTk�mg=F��m<mv���/=<s�HR�r�/h"�U4�����Z`�%[�R{���K	�6�4>	R����Ӑ���7�k��WT@���3�֗]G�m������w��Xu�c��T��^��oh<���7����䔤�OBb�c6�g"h�	@�(�R~]��?���b�ޞ�4��s�����4���O���I|�����*(~/����ޞDotS��q$mP�5X�^�	� ��V�8��C�"�9��wn��Ќ�
��b�=�LX���<�SW��[i�mo𗮤9�	�[�Ě\1ecO��0������~�3�0�C��x��%�.��r&)-�p�ނ�#{��@�P��*>#B%�B�����3�4�>1�MR��}:��W�Z�-<]0�ew����(=a~��d��������F��QI�u2<ъ�w����)�ᡐ�⠳����5CX|Z�sp��y��)����6��X7T�,�q�q�G]���TY½�+N��[�V��O@���\ y��?�.Od<4k2J����tғ$U�nc�TZ�	���?#�BTw<l\<8خ��tۭ��Yk�ɳ����ۨ5�g]PlQ닺��W��XW�˒K<�ޝ���[��s����M����k<��R꽊�+�S�f�����FZN���К��;��kB9d� �I!�e�fj�i�]-h{�6����T�ǣ��b�n�����8n0%���]B��+p��\K��)��H�p�8a�\^�~�9f
�AC����cU���!��VK4����� ���H��{����-��n����ֈo��p��I�e�؞1��R	��e��_��-^-?�_L�!R���%�Cj`Z���O|�A1�aK� �K:��4�e�kݔ���T�T)~��[6��Ҥu��V&���CP��A�g���+NNR�����3�N���=����BU��	��{�K�";�,K����[��vS�,���k!<'G��@��,V ^GtR�ïf{�m��dk���@a+�/��?U|t��&�	:N+��X��P�Koh~���˧fH�T4K��0��v��L`:�&5���&�T�vصL�CyhJ��$�2t�%���O�]��=mlu�o�y�G�z�32d75�>��Ϻ��3��Yp��VM�:/�	-�� Ɉ����zS
��u3�y2Dپ�+��� �VC�'"� (V�����i�����{���H�K�Gݺ�p�����K�_"s��:Քz�˧~я����C�Srsx�š$e��Ж�z|��hXr���R�0L+tbX�$�v�o�1�r!�5����T>>@߰'��/�����g�; k7�w9晱����7�|�^�dٵ�ƔX�e����y>]�e��+�n�/���ȭ`�I<b�g���l���y3��J_4G�$^,�9�Z ���w��Vw+?ccE�h��G��g��

}�n2�3=�a�������T�s"D|�Nzш"U����C�� �\tY��iv�,#��-�����i9�W���$�f,���B����u�N�9��R���/�H�J�X���k�S/��ͭ& ��$�6?��d�0*�!��j��{� ��)�v%��C~��|B�򱧏��'�v$���G�yȏd+�T�5kJ�	���G��H�m(D�|䉸�~l����m��S0��]�R�d��T� �>T阑��M=�4�@9�r�ݞ�U���H��4`Z�?w�N�^��{�ó�o>�P^	P�=�h��5�s��\���rt�b@^l�C[��V%������||qA�w���R�����i ����D��"��J)9_�շ�®~"^R��{�$|��	.��2�	�=�3����r�#b6�N�.^����>�F�J�z/� |����b�Zuv�&	�h'��y�d?�Htƙ��_X�� ��ՍN��Ȟ��#2��p�w`���e�;�\�vf���2]�z*m��6�O#�\��(>�C)t�oU��;�H��/t	X)Ѥ����a���w�?�.�4��IϹ�۝������
��O
8�8�#�u�e~�`�	`� xj�/���]B��I_q:�"zz��LL�
�{!mиͰ��+�0l�km�;��m�����;kT�@��'�!��7t��ɘ@�������8Y��g*J�aKK	�!0�%�K�P/�(�&z<ו%�~M�����*���.��"�gPǀw�]��Gxw^J��]�[�N `��wy�h��,',&ϨItr	� ��bh(%k���杊�j�=��9���\;�5��y�9~I8�����K׭Ȧ�$�'o�G��';=�S1��N�������R��l!X�lA�M�x��p��C�"���I5L>�u�����B��L%Z�	�۾�8��C�.N>��:�*/Q��e]gp�r/�r�U6w�%��!#J�@,���Iģ��)��2F��y�\%Մ 7{ ��
6�g��k� X#��]BFiXE�W��&g/��.��*+�ʪ_�����c��<xj�W�p��3Vm��S��߾t�����:���Hf�G�d\t���_eN��k���e�`�|J�>��Z��j��C#0�<&�[ۖH�����`FX3ΝE���C2I%��]�Lm�cߝ�!\�|vT�+��q�o��)�����f҄�n`Jr���ȝ�΀�s�h��8ԼLnk{�E�2п��-���G1�{�¤����{�|E�{��˾=,-�I���z�'���@���6����5��9V��UA��F�4L��Ң���܄������s|�z�RO}�P�t�8P�m6�[5+������H���C����������e\��z�?���+���ŏ᫏ /Ym�� W��q���q��T|<zr�Xhʫ,���{,<7�/9�{�{��sTʠ�:5g���N��H�}��g�!��}���K$�Þ�~�T�������M�v���^�#��X��� �n=����-��0�tSY�\Z`��/f��o���Dw����8�3噩Ȉn���YѦ;���$�P�WVH�	�O8#��:���3��y
˰��0՘�ۓ��M�#Ը���˪�p�Dd�.��O�±�$����.2)G)�/Z~V'