��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N'�|Z_&i��������GW%�12x
|�9�dΜ-7hj2k�wov�Ķٞ鳃�ͨ#`�y���>�P��Ac�=C:2�mt�+��Ɨg\��2O�|Y��Y�	4�Ae�+�}�U��M�:�t�<ؠ��:��)v�Ū��8�^�}��L�S�<f�%�x9d�1�����ԓF��CX����v��K�va���Q���	@�� ^"k�l�v*	 �b��)o�#2S�BŝW��B)����+�@f��@Lu�ZHb�)���6�'�y��z�r���h��Y����$�`�ˤ�)��L������<���s�n|���,��I9<G|�/�7�)/�r����`��D{z�c��Y���Eҁ�5���`eY�^������v��4g� c\�!��8�]�N�D���3(?yӎb��d�l�:�C��}
굑"��J�ڡ�h��[]c196���y�	u�բ�C��<6R�/����� ��k`f�����$�=��q�^��B�ם�l�(%�4�|>m/�.d��[k��9���U8�� �p�4(hQ�؋F=������Ov�/$e�a�����[3@������R�Q������Vs���	�ʈ�$mHr�"��x�<Xm8h���U����@|@�<5��'���r0�;���dBc���,טtu�H��1&���o��	��&�kº_+�	H;��#�϶�@�vd���],����h�plV�z����~�����u
`��;H�qM��{�4_+�0{�>d���{�`��	�&��X��A�/�|�e�TxgH���Ī̀#��I�^4G�NLj�ə<s��暌�<�͌$ja����*Ē���Է�T0Q����]�'{|4k��^RRV7AЯ�5�Hg�Yħ���8�y�����p�:[���i܅����3���ᡡ�v��R}��+�D. ���08S�]�0��fG��"T�U��E��IP�9�a�Q�U%,<�J�7N�P�/?O2�m7�����^۲�������0��fg�D��c��ftG��� ��W�b��n���)MD 3C�_^���]O�8��Z"1�W��2���G�Bs�П�!h���[TA�����/�X��@1.]ZV_��(�F�!�@�ߦ��H�2v;<UA�^oܖ�D��k��1X,u�I��q)'YӼPL�Å��X��7�ݞ����a��=�u�-�� ��ǌ�x�T�ue|���!?q+��k0@-XĿ���o��y����`>�y�o_*٧.o(#4AQ�|ľ��Pd4���T=J�Df�G�?�u����𻑤bʢ]��PY3��쿚�I�MX�\����
��6��e�	�zd(s����<*�g�ml�Hj��O��esf�g~M����@ԳZ�����3�`uC^�G�`��Ѩ'���5WdΓp0P@)�2?��^��E#N��� )D̳J1�r�,3���D�����9�Hc��I�z�ԏPR�S�zőv��]�(_��ó�U$�˧�%{��`�������
�0�fެ�M��J|�T"˼T�&A��Ӊ��R��*���y�iP����77����W��F�0�&X2�����I�����{�I�&��7�B��`LY�2k����+C�^D�y��+��٢# (���Z|�C��
;c���ౠ��L��t�s�)�=��b����2Sh�[*��o��9�x�s��k��RkYJ	ЙzB&���t�i=��P��~�f��*u.��=c�-ޏ��葜�O7�p#�рdQw�f��n��1�*���c�۬�YFl���浞��h4���R��}4���9��YK,�#����������L���+BCM|���?��<C!��f�w�Fh���D�8P=u��0uG�W�5�8<���c^���
��U����>�*�R��8�R�%����7��"���N�~���5�ߞ���r�_F	��Rp$�Ӯ�a��=�L�OU-u���$���=��?91�AM;#�a�{�I�"���477��e��V�o�B��X�m����K�E �V������T8�(�U�Op���WdUö�ԃ�g|�P5�u	v<�RQM~��޴�z��w-��Xy�d[�I��=z�q�޼��1�v��/R=y�>JAD��g�f��lb8=�Ż)�C�B��WpM�}�E��b4̼PF��"�!po~�|�^� 9�NA�O�$�
���s�Ԑfl��V�C(Q��e����IG������b8?���`}I��δ�{l~�����.(���VӮ����=��-w	�T]"�04
���e��k��@�3eO5�4]���d	'��8�|�eoȍ�vs1�`�R�I�r\pH]��K���E$@]׹�w�d�������O[ֳ<s���?E�	�۞�8Ç�x���N�Φ����>��R�2��ŗA�C�=����k~|��2�Q͇�J�p�ٺ�"�؁�V�3ck:bbHR3!�ӦA5��&Ea�:�)��&I�#�V^���>b.�/���.G��t����fؔ��Z���'�[9�HZ@9W��S��k�ӧ��Ac�6�W�s�&�Fp�<
����4ѼA��_L�����pQ�P%�EK�a�~�΋�#�w��Mu����I�q>�M�{�&I��<��̘�FE����t�?���I ��}�����E�s���Ţ(�?|A��ܠU�u��"��e�.D�b���CB�u��4쮗M���S�v��r�%�"�3�����+��=�ݖ����o_mDA�K�s@���7����^�ԏ (�+�\`t��N�Ce�*1��:^��mm�����b[o\h'
�S5T]�`&�0FGf�� � P��?�FƮG�Or]�� T�KJT�j��m�,�l+/���߾�H$����׬�`����]@�[+[�Q��`�Y�܌^�W�d@��-(Zw�O��O⟀���^����Qg��h[�}%��f���,���'t�	+�{�+s�m�dXX���^�`
�?j�M1���֐7l�>�p�e��6,G!��,��_����b���S�J�Q4��s������o������J�*�#��۹.��ouQ�ػ>ɾD�"��u��{�J���9��4�p�
�N۩�NYů�2��Gb�/�T��m���ţ�`>1	~��������]W����V��awؚGv�r�\�7V�b�n�޺)�^�f��s��ړF6B���q�?:�p����u��y�n�ر�Lۏ3�G&��f��O���/��}��Fٰ�CoD��R)E��:-[� �@'��KY�
A*u��9V>��~�8e�%f���5^�Ԍ�^��6�k}��;��`$�U�Ѹ�?-�����wQ�OXVN��ӨY�����V��{Un#�q�*<�,����&�0��r�>9����Xo��Ń!� ���,��Gj�䌠'������}WS:Y�-&$�/��S��c�&�8��"�xvk���n᠙|�T���ZJ_�g��0�q��D'��w|b�U��$`x�ھ?�zX�0E��U���áJJ��.��㍶Jw<�yV��Km�{	��_F���Ԩ2��c� !�m�pR��b�w���w`�"�����$s�G�����L���� EGw$X��G�(��[����%��0���OF�3QK�@�5ŧ��5)����|�DӞ�\�[�M��)+َ�����%�@t�qG"V�r}#�� ��;A�f�+1x6������Ǖ���/��������ܴoM'�`|���:Kݭ�Fc�B�1B�7�j
��
�m���j��u�W-
�6 d>�6�J��F֛T�3��22[�#�&����H��������_B������P��w�`5�8o�J�[�'򜼔�iK�ͯ���Zs(��&�žq-��|�[6�����$.��)�H��ص������4~�0��)? �ap�y��Y��;���� ��5�&�Fwbe���꧰з&�L��y�5X]��m&��$�}C�5�.�O/w�ʽ4�i��Z����J�=��c��L��ÐXFN�ުw͠�C�AW�P���Z\��\�`�|+硫���#sD�8�jbr�0ˆk�x��%=+cy�]�N_h+Ʈ�ca���O�*j7�Ӷ|�{xH��U�W�4L.QռMy[�xP���c���/j<x�uw�z�Pxӗ��RUl�~�NJV��]�D���͒������K9P��|?���UU&�fM�yC�0T�7�yJ�η=�1�Ot��[¿L�؂3��+,o*�q�[`o;4�>�B���R�T��qA�]7`�6E��5�ȝ:	�{G�]�r2J���2r_��H�~���M����Q�0�*<���S�-s{��gS����A�r�L�i=?7I� ��0ؙ�8�A�q�f{��<Z�Hh��.R�9ɗ��l�`��I�hc��!�=<�r���-'�W�b՞��pJ����j3���T���ى=��]{��W��n��5\����V��`=K% ��&ҕI�\��f��sA<�}��Al�1y�TZ��1�Z�h�Py���YGZ!ua�����A��&,Z�yN�+����D��)�`�� �y���'��ܗF�Ո�M�i������{g��߫)��U��s��60U0q�@�.q����V��'B�y�9r����}0�̫A'9�&RO0$��	R�Š��0�ƛ��<,��8�G��c��d\�I����,�{�2�h��Rg�+Hsȶ,���wr%��3���aGez������Wꍽұ)��b�^��\�ތXM>�������a5凥���-�2o�q=U�6-����/�~t�U�&��A3a���lkx3fhFg�	��
ߣՅ���oRvFmS�����	���#�����A�..O��8�ih-@Zm���{�&YyX�N{8���5���*�Z��[:*��T�N˗: ��(��١� J�<�hC���Hc�W�\'�����W��i�n�;�<!o�	A@�\��]A��j�Dm�!�UY.�"�&wޒ;u���/+�=W����m=�h�{�֤�2�x����ֽvGq��=MI�R�W�SE>ކyr`w�Q�D9=��9}�GN�%�;�j<`�gMVN��$\P>��H����8�LY_�X�z՞�fq�x�ŪӰޅS�k����a��$4<X"Hg�K2漷�e@w�R�u��tژ�1*1��V������eCT%�1������uh�1��f"F$�9����=އ?��c�OW�7�8$7�
�1o��_�`_9r��.d���D<�W1�ń��q|k��%����w/-9�Y:(vh'�q�ۙ�5�S�B�j�i�@~�=�:�
t2�&�B��酈}�KTe����8��d�\Z_���p��B�a�|~�����d��~B�����_E��5�zB\�l�~��c6�)~���
�%�'�f����h�7:���g*ʋ0�$��ɲ>iz�s��]�� �JI$H ��B0F1�!N��3@c�]4��Ȥ�'��5�$�x� c~�_�U�V4�� `�t/2�|�F8�b�9�a��k��prf;s�.��W�jI-e�!�˩2��uհy�������F���g5�؄}��]���6�ֵn��	M�z���!�C�Z��
l�̰��l�=�S�
�����֣^�lI9�(/p����y
����}ԐQ0ௐًoZk3ƈ�Hc�n^�)D�˺P&��@�w��J���z
��[e�,�~���`�Z�Xh�r7�h>�4�_��tl"���K� ���ɞk�z!C��i4F�G�n&#�z����v�q���j�ۉ����I24�_xB)��y�qG$7��W\[��X�q�!���a����~����ڌ���s���]1te�f���ˠ�f�/��@BR�U�p�fd\�D�4�jb��:o0��}�������/�`�b��O�}8�Yf�/�[����m��<>��++�O��*��L��`�Na��L����վOm�%~�?mX�ﲠ͓W& ���f���n�� R�۱Տ^��J�:�LLgd�K��y)'�q0�@�C�|d�іq�I����a��e���r��$�u���2���?Q�z�i_��W�V"�O�U��G������������ʡ�% ����e
/��ݵ�v����~�(�(�G�[8� ۫��j�;�Ғ#��Z'T�_W[['��/��Ӈ��(������Ң<H�n.��R��t�=����|�lm?9>C�6�(�����X�������nj�O�_�,]k�R�7j�;
�����^�b�m8b�T?Qs����v;�4Y���Z���j�����'[��B�T|��z)�D���ZC\=�E��r+i� ��������>|�����Y�6�\k;g�����đ³2�(W��g�o�>k�u0��uF��ut���S\l�}��+Jk����Q��)l�x��5M���k�7�㕠�?����k*�2�8^%տ}
Q�(��e�IS�T+"3��ʁwS�۲�;��w!C@��S���&�Վ7�|t�%�T̩��mj��~����<�W�(��HD���7*D�_I��z��@9Rp#���L���~E4,�R�w5o��굨��u��%S�W�p�E�I����^Gۛ����ׄ���师�͚VG���x�j�O����=m�X{|.�]W�������
G�w���}sw�����������&
/��������e�I�Z;Y0��z��U�V�Y$�se�&]���i���\+��Ew:�g��6������wn9�l�VO��7ON���,���Fw{�	
��ڛϠj��jG�ͺ�~Dx������k�kϮ��t1Q�#�J���g*(Yw�k;g;p��i���� �ە�LR�����wbuQm�}%�[_����W&�k5��4��Y�^�d5e�AL�8QC�D����U��T6L?�l�Z�N�}���l�'�$���z���ߔu(@���o�X|�{*��5V/�cn��B��#�ul�%�,d����������9>�|.x�q���������0����������Hi����U/�(�j0?���X�B�.{�I�_��@�;��?�Z�wCdߠ]4�h��t�pX������e
邏ߦւ�]e��6+2U֦����>=�&�y�Tk�v�Z�2bn�.����3.���9��j���<P�#knŜ6���9D$���\���������4��71�8GL����QL��*���W;/�7��͆�@	�j��=�w�\�LY��L,VdN��������"̵f+i��N9I�CuGj��0�b�C�{�v�������J���L�<f�Y�Oś�hH�l�t�c��~N�1�����e�s8������31�/�sr���6��y �&d'���͍�_W�Qï��[F/��oH͂��!������}��"�}���l�kҧ�8�q�*`�j��L9�����l`�{��>�Q�׶�,}1GWV�#�5HhH��n+D1"�S�ԗ��+��&|�܍��&"��<��7o�[!�j~^�n+�i`���>I���.���	D"��g�F�l�Zl�N������?��?��B>�d�`TD�6N��gz�-l_��x��'���,��eޛ��9��R����Ed��?x%y4�������x�
�٪I
���<�e��if\~��ռ[{�T�d�K*�G�U��&�o�"S��rI�%N��ǏSč%�����;,�*W��&�ZE0D�M�`16��\u{�z�YdBaPG�<�0G@���KÌ��{�,�8X�[����̜��-!��a&G�ˬ�s9~06ȅ%���>�.B�V2���BZ��"5tY`��3>�n�_VF�a�.�-w�ݞT.� 	b�}w� �ڤQd�"�4{�~I�yE2E���L��G$s���'�ߕ�̏yo�ʾt����+��hF����fzY���A�Ҳxq�G*��z�!鶲I2H�a��,.��2��#9�`�5N��O=�oː5�߁u�����o�����%P�.��d�� ��X��^_Bm3�5H~jx�.�\�j񞒅\�.�d�� ���pSP�|;XQ���i�~�녥g�3��nh̽� ��@�掬5_qT|.�%�3r��o��Д�����V楰�+@����ٳɅR��
u�`y]���y���7� nu		��l����K��\�xkAb09�W���k��܋K��bW�9�z5B�M�#y�siEF���?���b����l2�B�Ea_�!�-�}�D���O����̀{h(ա�{��)(���k�A�����O�?�b@�M+)�8Y}*:$!�
�D�!v� M��w�I�/J��J���II�em�:	=�K�����v��Yg��ul��e��?���h��[�*��l��l%���=pñMѕ��Nls���f�B��Md��g�2�	N*	�]��g�fylPc��Y
� ��|)��I'�d_u��
o�W�ݡ`�-��V7�#S)��b,^�aW����%��Q�����mi��l��:�͔��멂��2]��R+J2�10Ԅ�� T�̲v9V"T�È;�N�n5ӷ�]�0����u��3|���P�ă�2�3��F>짹�-egQj��fm���d���^}Td'v�(��A��15�?��0E^�y�>�lg�5h7HGԲ������Xl��,�U����-E޼|���[�YO,�bP��X���h��ּ[թ:������nG���ϧ�b��x�`g77�U,��w�Mt}��Y��Y�!뾳<Og�Ys�S�2�rg2�+Zݰ8*m]�+��6}�TS屃mP������C�:�.O�)��� Hš�{��x!K�2͹�]��h U£����'�hT����LSm���\�d�B�K���4.�'I���8�|�B�-_Yq<�MףE~=V��:��#b-�6��6)|���R�iK��7�ȭ?��.4�����G�r�����9ٖoL:V'�X1P�V&�~��$���莇��X��PIi��iF*#Z��3Jw]��������Zau�0F�������;���;��S�o]O�f�8�(`��	� ��ҿ\��/�&�¶� {:+��eo��~�yRE����s���rD�%��J�7�vMƗI^P��s���VG�\o�(tr���o(�qS�[lo�is���
Ο?)���i�سx��v3�-V�?���TJͅ�]��c����Д�jv����V����E� 0�$�����jP���ҴC3Z�����|�/��ʹ~�j�����O}E��ݴ�9S����kh�qB��$v��"��9��h����,;�����m�F �*=KwYf����/������r��:���G�]4���~~7-� ����a����sq����:�mKB�5Xm2W�38$�_I������J�X�
�_r��p^O��l+[:��z(�7̤���N��)�ߟY���Ǫ\���:%��eP�t��F7��F5B`@��9o#b�H�<f�F��Ѵ�{R܄���s���K�?��: x3��2�8�I┇��̟��oI�@W_��%剢������ā�Z�t������%WX2����k��q#K���:�F��� ��e3�_(�T�^8�y9aL'��h�L��8�[*g�ǻW�� 8�R
��E|u!�:D0\�i
�9��N�����A+�����ԇM�%"����cL0|���+3&���/w ���"AkU�a}"��N�sp���3|�8�ט+�!��Pqqޏ1'y�c�/�.�Ӻ�9;�Y�����t�/�а��x+�dt��=>�9���H�߳����q��d;���C���������`���0.Y���m�B�Oƺ�$���+zU����Ё��f�p�
�������ۇq���Ȧ�]ń>����;K=Cn*Y��3�(���xO����D7K����[pAnY'�Ż?����<��b����CW�v|үMRHl��4x-�A�H���#�h{>��P���{�-�a���'�l�V�C��س�_U�t6�4�3�	KV�՝R��"D�t���e5��T`N
g@��Z-��A���U=��r�%�ZX����ES1HH�X��F
�Rm�O���@y\���E7�<e�7�q�V/�����(ŗ��+�u޷9D�r�U��ܭ� �NO���wue�}����-�:���[@�!C��+!|���VÁ�ћ��c=<�5������T�L`�����T���m�w;)��I!
Ǖ�l˷����Ul��͖�OB��Ja�[�����,�bl8q��"�0��0|ݦf�}0~N@�Y��t��(�,c����>�J�2�>���\w�n�Sx�	;Aq�b�㞙W�j�L�c8��Os"W/�$C_����(�	�f�!E��e��y����Z�Ux�*���,�Bă�a\����9���D�6����K��Gа�Ϋqk�b>�J����7���Pq�]���&L>)q�-D��@����ɪR{�0o��>h��+����rD���1�p��Wm���6�k9���d�H�w�	�2;x�nm&8<&F��X�p,�������Ŏ������\&N*��3 x�B�{
#�z���l�@!�g5S�'+hAʘ#؅jϥ'x�cl~��Bev������4�֙�O��ݭmi]��AN�z����N����9�K��^�3I�4ֲÏ`7���M���%�!��N�sּ�T)Y��U!�9{?��	}O�kxD��ݝOQ;5����?��)�"�1���{��/�bU�X9�/����P�� ��m� {b{B��?�>v��ȇ7��kpNf;Ix$8Q��\�3�|+�(`I�P���ҳ����DcW�z�@�����J�����v7�6��S��+�o	!"1�Uf��,8���*�`
Ö ��c2��RD��]���z�rh�����*iC��>��V�a�����L(�����Λ����n\��Q�5H����L-b�Z�8%��<�~yX%н-}\����H@m��;�$�f%�_��&�Ӿ�y�;��6)R�!�,H�1�(��z5e���=S����4�-�B}�E�q1�D�@�2K9�ĒPo�Cs�\�� 2�h#Ҋ���C:r�i������-,`����߷��hHn`S�ϗg�ktPV��/��3'�����Uy��A°5hF<4��g�QG������$�x�k?�2m���(%�V>ж�x"(U"�(�K/��E�40�l�MV��+�)�Qk��쥢0٬�g����,�J����F��QLfK���r���e�d�8��a����9�J���8�'�˼d��;��;\�ېa׮GP�Z��U��lP~�@�D<@�u0u���<n��8��]�˧yG�g�Cϐ��Bm6X������lm4�$9�3��"�@�t�f�^ɭ��f��p����0�k?rۖ��-(��LKxv�/����O��Z7^&U5z����m�i�0�ؿ��"oq��ga}|2� L_B��9��E@
���8�2j�=hJN
��o'iֵ�5�wfDh������@�Ƭ-Vnض!�\p�k��+rҟ�p�b�-��ǰ�7YtԎ5�T㺤�8�������T���2���q��>�
&��Pᡁ�x�2�9��l{�Z)�rչ��4ʷ�+�'�<_����a3�7���::��':0�Wϋ +޿�Xd���o���U�M�K���"�|�l�RIV�V���Ȗ�Kkein�Bp�y��6�ycx��7� ����.�ù�Bw��Vz�@��d*�-&^x����םe�<��[(}E_�,�^��{6bD�%�&�^Y]Q��<A�8�WM���dj>8��g����t�0���L�����aW�(=�K%��Q��1�KKe`fF��u�z�./z� �����S��3����5 ٨��')��"\��'�m�xl�c髤L��J�K{�Z���l�F<�DI���$��{DK-�'��.�S9�ЂP�`Ӳ��Ϫ�4��T�/p|	�a��@�2��;�ZZ�����;]9�ȥ�t�d��+.dK,y��-���]�6��ʯ���q�]�k*)ɥ:��9A����[b��$1#Š;����'.�9�)��G@��")o�Y���-�ƭ�|G��;&���]��g]/ɘ�ue�y�b��O���?�j��_鉉�|�����V):��X|�$��;�U�K���Hd�h{ �L��zn�6PO=4]�O�iW�~�ܰ[W4�Ւ��P����Ѩ�Q�삅^f��E���l?�����f�u1�0���6�i��z#{b�x�݁H���B�aT$��]I�3r�L�;u-ǷG�NÑ@�����oF��h$�M��n����mM�1�{۷�b>��S�?����z������%���f�O�}�o���Z׻���QK�[�'��Q��9�P��E��'Ux���0<fAǰH��}�#�́'�~�#�+c�4#bd8<��s������}o@��LAa�Bb��N�+�n�y�ęI��$�
��tI�U`3�vֳ��C$�h��p@��]֜��k�Υ�0~'x��]&~ŕ�]O�M���\�@y��(m�	�ʮ�Ք���o6@����#>z<��� Y���@z�P�Bc�-E=H������7�I���bX�M��NX_�>�&��|_F/͏_mR�U��uRK�<��׌��������'0���IlG#����,	��B�����WK^&��LCՈFC �#�霊��O	�<T5~�����nk-5�Xw7|��e�R�ǹ��̯u�k���cњ�5�|�Cs���=h�y��v���J�m�ـB�a'pd�3NU(�9i�TM�-iVX�rS�3*���οR��znN)PQ�Y�g )�>�UL��Nb�	��ՠ�k���D����m�Zv�^�q��{���� ����)�4��u���w������JQO$fF�<�ΪK��$�{~%����E���0[��f�P�khC� ������U�<$.��۱4�Y)��ɉ�X����N#؋-��:��w�pyR�2����A�&v<�S�?rw��@~	�Ks0d+*0��5����Ŀ"N��GO"t3��q�
G��ڂT�Ɔ����\'m�/l�waxa�g��F���I�*o��%��#xF���%��u2lǔ� F�/�����BHL��Ā=g=+�lh�RB�Nֽ"+��KÍH��,� ^\Č��o���ڽ����x�#���8���A�� �z��؃
�]Җ.���ɕ�Lg�m쮂&-��))�F���Ұq���89���/|�8p���0�n������b�:42����ɩ���8f����̑d�L��~ҾK#B�׷�ה��_ڋ?X<��n<y�V�*��e W�)�]���b5��� 3�M��1��뭋7���.�v%"2���YWĬj0{��˓"�YD�IuD�Q恡��at��*0������!qNGD]�#���c���2��g�'I������=��j��CF'y�kt����K�����@�N���x�:�p�?� �fkD�V��	��bR���%Kت��F�v�zNd�����҂=�>��kA?��A�V�M���EJH��˸��G�uj�ȡ�	��J�F�f�W=Ÿλl�m�$f�vڄ<�H��6�J�Hӡ��R�k�K�hZ�%�\�I��%�ָ�L��"��-RϺ�]�<n�3��9���.]�܄Qܵ먔��� K���W`f���_Ռ؏�	��e���d�������^�.G[̯��N�)�+���>s^
R��E��=sZG?��h�7���0�|r���l2N&����aɷu�H�� ����w�}<)YsD$s�A6�)�����U���Lm��\v����"��#ki���z�I��pL��]t�����;�@����o=�j����N���ˢb>��`U�6a�y2/�'�+.v�x��?��Xw�5��p��c�p�/����4I�/�E�����<a&ř3��b@R�c}at(�s4Fas7Gڲ�k�2�������_v^�g/i�:����N"M���$�X�\��J�HR�oj�#��P�t�#����1��/�r������߀�����V�ߐ
G�����iXf��s��� ���;����q0�$�c��?�����t���r]k0y���+?��k��:������<�`OUa�^��zBzN�T ��މlG��`$cnu���.p�dU�6f�&�>G������]��H��$���*�Jͣ�h8���s����9yX B!�.��W�~��04��2f ��E�,��!�J�(�	@A�>�"ƑX��I�����K���E�����!���q��3�`硼�A[.[/��o�� Vkq�հJ��n���L����s�Nֽ{�>�<HRυ;����A�&2J�:.ϔ��=n�Byp�P�­�nx�%�:	��l1s9?�ѕ/��� 6��&AL�Q�c�C����r��%sOg�a�c�����
;ta0CL��}/&���=�ۑp��!��ȣ�����๧�IY8š��!�������8��Bߍk�8Z��]|��p�Pq�P�'#�M���'P��P���D K��q��"ŏ��+p�k��D�.5����&X(�41�fH���k�>��=���N��
f`��~ݐĳ�����8olۼ��Q�h�Q��#p��:�*r/��a:w�(�TG΃���|~#ŽM�j�P�r��`��Z~�mϾ8 }�b@C+�h���^���j���f:�	�{7pr��v��k�m����{j��S~ւ�+j�mM&r����C�^�U�:(����G#*z����7��fAӡy��p�����Z>�Op�ɪ�&Uo�\'�������������1�;�L�)t��I���F�R�^JY�H�&��+�Ԋ{��ߛb��e���>P�#l�C%�B���hk9v�!O�zq�x�a�cE��r��=ۤL���>((\4a�}�Mm�dK������֯��I,�_|�� �6��I��aF�n��HtZ��esOy!��g�}����r��R�q�$x���Hu��FE�R�$�ne�N�l�%�O�id�}�q�/�7OJ��R��V���_q�Y�#T�羜uoR����M֮P����s�y��������H�s�}K���f�Bw͔@�U��2ߣ,^z�] ���)!ɻ�,7 =�W'.=���6KEĺ8��`_� #i�@�C"�2P���B2���Ü������f�^	�m�q�5��<vçQ���S=�:�-3��)d<�s�U�JU�I�{�� J�b��'�U8��`:�#O�3��ͼ��{��dp�E�Z�F@ɜP+I�	ȵ��8�4S�f���tq�*$���*�\~����@��$��/$Ͽ�ل�Z�H8�Z�I���|�z5�i���A`tZ�ٻe���
�k���hү	6�ͦD4n�4�1!�TaÍ���.9)�+�������<�sr������uQ6#�c��B��5��:Ű����zB���:0�[G���ÿX�w�	�������R�������W� �r�0�sc��F����:��yI�7N�f;���i��p䷏��.��]�꺩X�8���<n`�ԥ�[�鉮�'�����`�h
�M�?�Z�h�a����&��Uke����(:��}7+����zR��@��;*�vN�H�A~b�����lW;/ ���$Db	�+�J�HGW٦�g�aq/��*��x=�DY��o�H��P�ҮЇnp'����L-Iut���\}i˯��g$�/��F�U
*�M�Q=^��
so|t��D}
)&/C
��u�4r��E�'��:i�^�����ō���z(�i�vlD��jˀ���
i^�S-6;��~���EK��?I�9��8n��?��P��:��H�~�Ĉ�4�(>��-���	!��# �m�?���~���5*��R	̨g4�8h[D���Hv��x�؞�U��0�����^t9�mW��GK	�b�֝/E��#䲍p��k��
�J鳇z8�?��V��P���d��:�*d+�G�UjuN������������r &��(�ة��~*H�pg��4�	�+�������K�c䒤t��n���5���	�Y��^���G��{�����g��4���FJ�j}�Z2�v�'��"p]8,�5��܈�H8��Jv<�a�a����L��������s�r�����O]�=�%�w;�	֥�]��P�l��U����Ѓ?��7x��
�.�u�-3x�6 ����.���f��%qڦUA5����~O�?W����X}k/�m�q_�4w=~E&�87���	�kq�X*����$�o�bzY�^4��kSi20��g6��Y�WG?	�Qg���\W�����( s'y�҉��v]0�9;_͊z�ֳ�]�2\-���&���5��t�B��xK�z����}h�гh���~o\>L�����
7,U˅�3z3��@Oɴ-���3� ���{K�
�y%�G�7��&��l}5N(io��z�Q�W��pe���d�����CS�!L�0m4z2�s�P�* �>1i����=�!����v�Z�[��jDB��$gV��y��i� baZ^D����N��^�ܢl���Q<�>��!��-W�6^w�������>o��zU��u�;G���+|��|����'�(��]������p����hA�fQD� ��{w;u��I&�S��d5{wt�n硾c�`q�B#速}�j\~�z2 	O��N26�ө�>�Z��W>U�=�h�ļ"�"zv���D�r���Uq�o�����_mq�ǽm�Yo�������q�2�jڐ��66DDϛ��������S: .U�Q<R��C�%��}e��;��f��ԣ���.]G_V�ȇl��d�8�c'�� ��L�2�%��E�Tb-�&CptxT)i�@��ۥa�����CW��Fz��������Mp!9�D�x�V�s��.�A�h[=�Z�6 �_a՜�i��/��X�����"e	���!���؆������78�R"w!��ב����hO�v�P�~ �ۄ�}r�W�,�eW������h(חm�2���+�n�i�ɛ��[}�R�t�.��Ԡ��sv�7�mn�*������Ҏ���
�̕��'B�T2��?��Nk�*�Iz�a����S?�S-ACQ��UR���n��@f��o�2td.�ϥwq�'����Z_��z�ᒞ���Җ���A�K�\z�U�Sb��%6J�{-��M�^���t�o�WU�uVdš�f��
=<�|���\�v���,���Z������Ҥ}�D9B�+�|���%�d�W�ӦQ8*�ȁ�'b���I�G[�U!\/�u�c�U�������63����|�jH��R-nN�k��Ph4�նdR��p-VƆ�&~�`����Q��Z����|��/��;���D��	u	��M{-�������������{%���^>� �I�˱�D[�Zۈ_f'�j��ّ�	z��S-��u��o+~d��]گ���,v.��>�Y��K�Zn��0L��{0k��5�K���3:�?����^�����k<[��/�ǡ 1M�๮��6h�d��[Zm�t��E{��7p��f���  :��u�ePl�NȊu̓�l�H�Gj��G1CIG��+n��Kn�$[ �6M�(�WY��VŉaL���}A�Pot2�7�у���W\A���e���\���a#�z�{��X�1�:LI��8x�@婊����g: >����*�o��Wg�=T\�2g�	2gf�����uT�LO�bЖ�k����15��'0J��{���˪p�>XZ�6r	�k�p��l_���DU3 �Ƙt�W��I��s?�l�pu�ƒyد?�4��7F�|�Fp�p_���}�Z
��q�O��F�˚�K44	��v[�+�y�w��=�ہ�Y�
.A�=�n���5\k�Fb�������<F���`�#O'�<�f&�s����4b
�N�Sѵmׄp*�:*<yz�5���u�"e����U�irU�Fkg�"2Z�D����m]	[]j֙<��\du���j'�2���⮭v��w�)�}��yns�m���FΩ����`7��FS����"��fY1+ۂ���3���n �R~��Gt-�s�;l-�fO�	���v���.ÄS��W�~}�;m�����89�:�Q���E��(���3�����f��l�� ޵p� Wt�P��8�4,=��i�Y@�i]*�W�� `�(8[���Pؙ�Q� �ܔ�QUX倹O�J�}��H+�B�>}�{e�d_k����e""�< }���dZN�Ǘ8����|���?�JVD}�e��qG[�Z+�^�x?-���Vҿ�f�~�����L��2��-U26U^GU��=>����ˇ��>�C�:�j�t_ϓ��㚡��������n�F�.i$�",E���e|�J���gmSN��s��v�o�6E:�r48�1�i�[�������@3���٪��/���cLRn�
.�
�A�嗁�x6�Ē���ysw��lv�=Dc��O[���Ƀ�8�����d�pP`'�J�I�����J�NHpaQ��oH�+������<76�>����!Q2� m~��x�#�C�)�˂��q!��r�I�oGDz�}�p�q%��d2S沆��Êq]��֣?q����R�ؖ�جl�k�<R���"|��X�K��OB`$�< �q�P�8uv pG�\b�2�6�h�m�	6��ZC��dv)�wZ �G�q�+�� �7J��Cv��/�a��#wWV��X�л�� ����AW'JN�����F��U)�H���"�^�C>��$=�����\z�O�SK���b�1U2�Fo�8����Yw�0�CYX��r���΂�Y8�<l���:1AB:�J��Y�<�����g|�?s�z]t���4N���P�uQ]�{߫qI/���(
1yX�ݾ�J�̂���D9�<ߥ�a�����EI1B�~҉�$�x
�ޚ��g}Ϫ��}���V��''�?q�pyʔ�@�z�}Ń�fn
{�Dh54�H m��b_�PzF��ǌ��H3��Qqt������:a�����4Q�1��mH�I���řh=����k0O���V�F(�5�C���đB�`�P����Ԃ����@#+N_�K4��k�����}��m���f�fhyr��YSu��h��2���T���x���8�)uST�c]Lk2U� a{���]�nVֳ6�6�Z����$U2�vQ�	ED��� 3,;)ֱ�Tj<R��&��,
M�kܑF�ꈔu�M+��ʴ?z� ��BҒ��e/-.�x�3��Jp��D�IKx%�s���F��H�Q�\�R2�dg=J���h��^p�YOj����e�P�l��9q��L��LI�xA7O\�9�����F�#�&]��Qwfį��y��y��!Y��Cm��,�Od�+���C`N�_F9�
�,_$3��d�x���6s���b̑Ij����!��.�E�@��R�ؿJ(�N3U�V���%�2�g�oxdN���пh���Z�L]%�v��WN�DX� :�o0�_�SQmp�d��;�:�?K�f���&oM[:��h�>Cl)���*�� R�j�rE�E
��]���_���|�$�V��t��X"M�w(�i��,��-u�o
��aϿ_hY\	��>s��Ę�����l2�o��9�%W(2�>��5�1x�^�-.a��YXѰ��Q�Ed��ˀ��}GH~���|,"ˎ� ���S�%���ťg��Q���w�4)T�W6�u��}*�QG��i��l�Ҡ[�M��n]��DN��@S�\���4��r(v4fU��覓B��}Uԣ�/C��d9C6M��]*��:愌���D��-Q3�M��X3&��(c�IR�S=T�Ō��w�*U��R�
;{�{.ƴ���-���4 )B?�Ւ����3FLo%��3��h;�V㒙�� &�g!��V�U���Ny��1o�3�+^Vp�F��9CR:?�Zת�`����t�2�����K%��B���Y��^�V��bcjs�������l���J!�]=��c�V�Y���>g���Rc@�Q�m��t�X�G�"
/,9���KYrވI��Ќ��oPK��Qʂe̙@�FzAG�˥X�Z]s��\�|��A�%��$���)&���ܤvvI�n�S�}��!�Z����݅�V�{���2�ޥ��~��P�zʲ��3�W2����sN2aw¼^�o\]���f����D�[T[����g|	�͝=We#W��D&�ՈZ��@��)$�&���u2������-$�?QO�M��|{�D<0���4H���h��|0�qHew~��_V��ۏ�͘������,Z-/�0���s�L��"k�h&U�m!�[��eEXf�3Ux�[�F�<���Ef��!{+���9��v?�,8��A�-*�Q5	�w�W�:��Vp��7F�5�n�-����J�~�멏������L�*�(��Z��d����N�!��X�@{H]�x�	.~�D}tk��?G%��W�,�n��2�x_�:��`H��aE�PUC
@���ɫ�)���m��*�2DS�M
�o���yRȋ�N�\W�T�RU���jh{<ƣ}�IdCd�r�e��vc]���_>q�M�0�}��x�QlЊ=oޟ-Ni38Q����sS���	}���'6�E�Θ��� ��)D8:��E"�44ӡ@�3ted��m�b�e���
ˑ�5G����)��Mi�k�����úv"9�Q;,����u��j�%+�k{d��{h���-�~|;�=��w�
-z1n�j/�垔�����>�e)u8^����O���/C����T��|]S�8�n�n��v@rV�A5@��RF-�y�c�>�c
~�Mis/�Gї��,i�-����K�Q|!%ZpT��iq&B
�A>m�b��V�x����m,�0�Fr�>HȀr�Jf{����:c�n�*|����~�����-��pv�E<R!�I���EG/t�gm��ϥ�L����i}Kdc���xD>�εq��j���4���R=���)�([�nФ9KF�_��y�B(����v��*)�g��?�u�A��N���cEj�I�/X���n����W�������
ez�	�@Y4G|�^t�y����'�6?_�So.��<u�i�i:_�>3����3j����O
_�96|�� �;F���M<T�r7��`3��)��#��:�����	�i��$���_����QH�p�� s�x�X�<Z�jUZ����x�Z?U�=4BڕY��9�S�칚=ê'�v�f��+�'|�t<�MC�(86u�3��	�S�C)߂�ئ�SB6G53oa�$���n6G5�QL�G�qD*p�k�x͇}'<S�@�'��z�Hb�d
ޫ�yͲ���|�ِ
ҕG�
c�ޣ�_"��s|��FbnȹDz`�����a�d#�'�`3c�^�
j~��nC�B&d*�6L4��a�|CU�Zg���[�PH ����|9���k�(ջ�^���&�Ns��@�[��4=yĔ��g}�՗^`��@#Y�w�&���|[	����s_+��!�H��E݄	���h%Q�<���Oe�����x�)�����::��
�6Q�J�.������Y�;�$���8
+uK���)D�8V�^5V%7�������NI��t�������Dk6��d6��F@���-�� !�q���� �.�/��;�#�.�C��ʆƛa�"��9u�'~�V��(�K��OU�u�R\0����es�}��0޲�'�O6|z �-���2-��;Y�~J�?�iӳ&	�KLdg�A�9\iYn�'�$3�4Ţ���W/O����U[[!��m<;/#�f��y���A��-�Ѿ5��V��|ү�@q��˦�GR����f�؈M;������5��ڱ,FF�]�D�/��6�1xN�����V���X	u������g�� .�t�H��a�[��;�ܿ�\�d>�4t@�%����Ԭ�#�,� �M�>j
d;��H�!�7 �]%Q־�t�a$��j����_et&�)�ñ�2(#U!t%�+��<67�u�q$�Z��2~��*�%��#��c�/��c7���6�EֹVk�Ϛ	�x��)o���p�������RWHd� �/�^�~�˅O>�.9cn�Eb�d�Cn�8$�;�J8�?�|��k\e۞��w��o*r\,�Vd��e*;�̱�*k
.�a�q�7�~LQ�T�SJ�U�&��AScv�Q�,��ӊҦ�d.��rH�U~��dN�flO4� �q}ت$�]�^G���wF�-�tM�N=�׫>a�˨T�%�?������~�v�'R������{�R�n#��T���8_� ���}���2��w쮬c�;+��>����T3��e,�M�N	����D�iՠ\�}�:gU�b���G\An=�K���1��gX� �t�
��ֆb�d�g���I��G YI^Q[ɋS����s���SjF��G��(��� �1�;�b'	v��y�	����7X����(���H��Y��|$��hP�`�+�eڞ�m�:�s��_io��,��ebX�E�%�w>�lI:���#('JZ���t`����Z�_	A��37�?�nx��G�����P�&^���&KUFWio1u|S C��^_Ns��|���Xf,'�֫os�v�mt5�S)?eS�)σ'͉;������f���'~��da27t.������3�;�'K����k8��e���c��4�T������IVl��!,��9�
p���_�-�G�F���6�lќ"ցZ�n���M�����:�7/ҵ`w����(|3��l�YUV�1��ׅ�Hh[�e�ꍆ�,\)F�K5�Y��	f; ���nl��<�O��$�:@��L��NN�<ŉ��ʞ�DNW���΋�8'�J��))�(|���M��*O�'"��u����ד�K;�x�F�|s!�V83����$z�q�ԡ��Í����ޟ��Q��$�E_XM�b~�#�u��ʻR���<�yr�0�W�$��$���"H��0ho�2e���4�n�c�N`�a8\�k2鰓�"�
E�}�A9]�H�F�a������ۺ1��9�?�i�'P�s6/g���fF)R��O�g�f�[�'���E��j��:���Mog�ǭ��*���= �Q���K������0�w��������Q�e-l��BR���p|���+��'>������+���w���O�,���>�&�=�ɪ��7qy�����3/��)qYJX�C�K�Z���ƴ6鐏��?��K���>����`�v������7Alƕ�@����ѳ���zp�,���v[�r]@��`Y�0����tŘ�����[a����>��	\����2o�����X�ֵp ��rXMs�7��J�@=�5���º1���!1&}09y �eyO1
a��^�/<p����H5�wT�=؊Z.
�\�އt��U�z�s[�L3�*{-v{�E����v�4I�,S�i�Q��eň7����^��s��+�9
����*./��;(���`lݜ��L<�8�� ڂ�Q�o��~��G� �)���@$�2!Z�����V̀ܓ��	�j/�n���\b�N���SJO��2w���e	�f��J<SgQ����P�I�]e2�R+Ffx��5RU�ޤ]�5��fr����1߮S"�RBe@� .��v!T{�G~�"�Mp������D�����R�U��Ce{H�����?51�v��b�lr?�4����C dI��hb�=����i8&�+h��4�S��:���Q��Q�כF����O&?K@�������xF�C���7�s�ѳ̢A�0��myq�~8Lx���:9ܛGwy�����b���Qn�(�СF�?y�݇ ��Q�M�NpW��p�嬚8d�6H4����CZ��3����H>����z�:fE��Yl�v�g���yS6,�$�F8Fqi���i��k�u�0E��w���q���Ҡ���b-�Jǫ�is��"�um�Y����U�v�S�\�i���g���+2>Z���n��`wz�R+@��d�������F�����ùRu^ۥ��w^ΙJn���?W��%��s��<sf;�C{��T?�5��,=�h���wޑ�>1Q@x���,�Ѧ��ǻ"r���r囈։��pGa�ц��l�w�H6O���n�s8�R�C|�����4X��
�RCt�8Va>
�噿�v:]A��8�ds�����yi�Ak���Ϭ�?:�9)w��E��s0�8��"�8�����[ �p�����mm��\bs������QZt
?�����@(E9�X�j΅�-9(d%,�e�C�����l^E����7�c�Je�
�{�@L�����kY�_a!��#� a�vdeL�u���-�UlB���~x����p3�cr��$GIqT貫�k�mGqF� ��bc{=P	gCܝȅ>���󙶔���!�z@s�P�F0��)�DRen��q-�p�so����z#�BD�
b�6�p:^����Nr�`4�{�T�hrV
��Ƞ�p��[5�@��(t9 �>,h�x����,�.6�B�_Ƴ���IӢߪ�8���WC��ӧY�����M�;��s*$v�	~hl�޺��*G($E���m�Զ��s��8�N��U���վ�K�X�*�������q���љfH��<� �A�/	 �](�Z^�����xZL�z��>� ��c��0�w/+�5�Ùu������&�f��s�a5n�oL�[.#R7�,sHw��*�*��#��ZOi�s�Q�;؂E)6�9�hs�ꔕ
�+?Hڜ��(<Z�M�%.L���2f�74����K�+�(26cK��7�j-������Ǎ��U$��s(_����~�Y ���O��Ag��S{w#�s����GO�x�:*Q^�?	֎iG�{�_���(L�4PA�w[���0Ҭk�e� I�,C�g^���� O����/9�r1yME�\�(͆����o9LS���Cᜨ�ظ�U�O&*>����y�=�mW� -b�'?��+�	��n%�Z`Ų�N�m,����:ٯ�#hF���X�MS`��& /qJ�5=�v0��/6����ɿN�JPԙ�~�.A!�)�n�J�$�Ĝ�[O��/�����	x7��,�&IT�>�Xp5�]�]���O�i!�G�@�;5 (�<�^b�SC�|[�'I��~#�^&tiI}���_{���9\�r�I�\�K�!w�IUu���nב���B$W�1�2��_�G�-g:�E�y��to���7��WP�Ki�5��f��۫��:Pq`�jw�H^�����)����A]TIk�ǂ��6��sA
�ZA��]}�e]�N!`ᙷ!RX5�9��^�SB�e���)���-4̦��Q��D}$Ց��9�_��p 5�Z!]��NB�v���E[x��*!s%��_==���n��;ħ�M]��%�+��΅��?ݷ�&����=R�Ua��"f%a֟�|�Z+=_ͼ��77{�~k�%"����:ٵިy�"�ɦ�"�>i�k�+N�IOoݍ�]HIJ�:N��ꌩ�������E�O`��[3�'��f0R�.ض߶���(SL��:'��pH�ǭ&��a%�m���=��0�(!؋3�I�ݷ��fn�X�u�daW�����%N�,�d��ѧi����W-�P��	�\��u��0(�ю)��8᝗L�坨Xq���'v�jD������ϴ.z�$�H��^���o0�yޣ��r�����ԃ<GԧǋD�(���<�B}���<�	P�����"Y.x���ZT��[Ä-�jYqG�9�ƙ�/;܁4��Z	�b+_h�TV�C�H���!m c*����H�`��ͳ@��&,yQ������u��# גT!�
�[N+ݡ|,
JĔ�s�S<WQ���T��9�C}��}'26�a�`8?6Q#b��F�_%�g8�Q�1R:�Cnw�S�]�� N��)��<��^��)�4>Nռ���v�(�e^Ӻ�ߌ�xad:j4�l��$�팮5zq��A�A�J2)�|,�s�������a����/��S2C���ֲ�39�;�[@G�Dͯc��(�*�Z�!�T��q�0���Ai3F��H4Cw�����H�|��-��r�����[H>W�۫A���c���eZ �a���l&r|Ǚ��ť��a �>���/!Rr��E�[h��䷅�t�����2���&c[0G��D?�������.��1��c�WM()�J�=�ɦ��Gp��w��Tb	�� �������s<I���g^�)�vJqN��� 냆w�E����P{��?\y�����ת8�e��Hv�ªlC�L]z�IFn�,��I���8�v�Bja�M�b������5�<����X
���P�E+�yV��,�휩�{Ut���w�6�B�j�`�+B�̓a1+����H4�n��:W��;³=�!��K0(��:"}2E�ԝ{��722����?�``Z��r�H�P�C��|�n:�נ�>���L�D��M$N��A�m���ކ(�LL�z����ؐ���;�D�=7҆J���+7� щ���/CF&s�ׯ��?�-uV�ӝ3yT�2�MB̉J �Ǔ��g�ϒ���;�F��ڭ�.�����q��S	VՔ?l$��r\>�]m���'��i[��#�5{n߲�Yl R4��&�j�u�5�E ߨ��s�0ɀ+��䂌�~<ܟv���~�����Or+e�[(�S~$�dr@Y�;���o��!7�N�w��gq�tqG����է��ޥ��N.0�zYГg�lQ��vԚ_��D�P*k�B'�C܏�{f��L5w�4����.4Q�'n�:���b���%��v8��6�{0��