��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��P��=:� ����(�)3�� 5����l]0�ك[�Y�qޡ�(���fZ��#b�}a�3�
>cO��o�LW��4�C���(C��&{��"�v11#/I�&�)�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)NU6�06�
aa�f�˥c�b�.hǣ�Q����9<���A����&�OGW&�NAP��~��K��#)_W"s	�q�w�����	��{�C�#kaA��Ǝ��_�,֧�H��N�ʨ"�k9(�V�}�HG;t~��jLTz�T1�����I��[͛�k"�dn�Ks$+� s9��wy�]��ښ~�K���uT�~&j
o�&;��ʤ�CC��'��I�?+�,V��Y�u�
���&ihfg�ۘ)qb������F$�.7��S� ���@|���I^������t�t����z,a����,�	`�M6?	�Ni"0K YJ>a�[�6�x�!s��X߶ș\.��Om��˰�뺧S�n����QXcF§P��x �
�8��8_a�
L��4�~���J�����u�#���E��3"M���Sަ�Wr��Ҝ�N��ʮ��ᰥ�K("qz��OQBx.�;���H`�ApR�nM�  �����Zj��z�N#~,[���n����VD �]`�A������)���L�������,�Q�b"��$��5
dgV�Q�7hHh.�3���.���RܒR�Qv�ҁ�0�û0��g���"w������5=�bTŇʹZ)�����NP�t��#��eMQΛ�)�)�)w��,�_Ӟ�SI���&����S��"���Q��n]���������lȾ�[�JT^�wo
Mk`fDf�b1�D4�JO:��#S�US��?	�JU���0���AQ$�k��K�(��&cOd���L)u���a�aH7u��w�A�a��&�O�cm�{����cf��'�,u���@_�J�%����w�';,�/�?�cN���ɶ�� O�	w�"��ib�}N
vl9��fK�����/�5�� ����G7&���>�)aq�Iԉn�g�w����e��{(K�~Lx��h�SjdX����l@�QA�-4Tm���f�@��
�*�'�;�W�P�VՉ��� 5����Ҍ�E���N$��8�V��������i���$N����ԕ+n`���%��Q��������v�;<���t*���o�F��U��l��KQB�^�c:��H�&�ձ2��Bb����\�'zH�:�L冓=+��;6��7	�V ��_Y[)>[����9{w��|q5(�؞���hW���G$w�S�e����W��W��dҾ$�ðd��hw.랙���Qn�[*���>���ݦ��x�H�t:h��Ҵ�R!�筎y�9��Uނ��*��2�^^;�n��5B:�X��1~�����w�1��#��]��;�@��j�^E�����h�;ʍ"���j:�Ú�F��)���|�gx����<�s��N�l���ܜ7QD	J#[L�3�T"d���3��ȍ�M��v�w@��� �}p B��s��}���{�q��\�W�IӨ�����~�e���y��\���7�OK>.]�$n8�}}|_(3>�&�<^��U4�.So�~8�no����	n���i��}�f�����a��I'�Si��"���|���G\~9���AH��sC �Q.�I�κ�햇�
�i�YrZ�DU��[1�c��uI	ڒd?�Tx��h��(��`�:O�j#0`���� Ԓ(��/,��62�
�(]
=<�v���*��`uա�=M�����{*p���1��-C�����&{��[߄�yȥ-�y�W�7:�w��#���ɑ�|�$M�o���$���4�o6$rQt�S�]�}���pN�#HY�˧�k@+m�0��K`^�Q���L<o�?���zm�V�#�ub�)���I�dX3��_��*S��_�G�h��Y����ר��$���ژ���c�F)Od�
�@k@��� r�:��i�F����̙�Ac���5� �*0�i����)х��d;(d|0a��r������ѣfTu���&��E�z ���>�=Lڋ�M{W?1U�	f�ִ�w"c^����l�E���d�g\G^�%Ad ��$� _�I�3�շӢ �����rnp�杤*�ug�@�US�&HރlW��I,6KJ4�z�_��3�?qa�Ա��� s����W}���}�+ �ʣ!Y������4Z���!ʑke��y��7ۡ��`��xԴ�l}���u.��P*���S,��o��~Q2＜��U4�`k,>���8��a����׷Z'^ˍI�D��<u!�Ħ�vH���娫W��b���4��'*�d�~.[I��D�:߰���$��\}�)����Sy�e7���K6��	T����>�z,�i,+�Ò�wn8�<Wc�Ի������ꃪ0d����m�|�{C�s��ᩀ�f�lp범N��X
.�a�iØݧ�Y��|��T�!�B�a�Qٌ̾m��O�d�= �7Qx� B�GE��w���([�R��wI2B��'Q��W�.��y	/5;�u'��^��a��:o��+�P��;����/uW�
����fTt���e�G�زH�A�k��Rηk=�dr�?b�d�x���+AjMk�F�|��U������{R�\�x�:
O��W�(������N *�az�b-눙����Wǔ՝���0x��a#��¥}�`�#�fy%��Kf�bLq�銐��80Nus�է�{8�~�)�L8(5ߑ"U�9���;��bN������~b�g�
�goJ1�`����z��� O�R��<�C���a��S�\���u?���-y}kLZ;;��Q��aɔ*k]�"ړ4c��-I������=l@k3̸w���T�K�3�fHb��~4?���n���..��.��n�H`���BY�����5��<�l��U��?���$a��~��LqR�M5Qu��p{���]y5/&W|����9��o�^��M���l��W�����R�����硺̖ivmIz�z.@��Y�r�$:�����Z#����\���?7��+_#�3�mj���#"�+�K����~MT�`�pT��vҡO5Is���Y0���^���
�� .�_�AU��4�3� �����g��ʹ)a?Wr�5�;�PR�kS~�s����5��3Q�PYNgg���5g�]5 �˿��kT}�9��NX�����{�2A��=@��?)��Ը���}"@B��H
�:�Lk\F����?�p�TM�A�u�_U%�Cj,&{'�*YF�+T�/�$i�,�����X�]j��b�}��G��s�]�nX������c�uX�0�q��·��t���k{�̼X�%@��SG��}��ժd8�:�H����"���1X�$�V���B���g�\�˂0)%w3	C�w��W� �����oW>�gZ����	: �݄�QR�)����n��A���5n�T��q����h>
.�e�{Ԟ��Ǫ�����η��r�>��e=84ݫ�M��rxȿ��������x���}�~�3I��ϳv�������a�߿���s�(���+sG��ZLօ+`{�Ǡb`L�5_���m�e�F�g@ڕ��5�~���,}x�n,�`�&��pڰ�A4�6�o+�����E8J�'�σ���G��v�[�����~�Vɏڨ::�ꨛ��o>���������N%�9�ّ�a�<x�y)��Шq���6�^�\��U'P	ZI>��M�}�<�l4�;������f����d�k����{/FY��>��/�hX��1Mj��׹E=*���Xh�D�E�Ԃ���Ӱ��L�{�'÷�u��7��bc�	�݆�D0�}�!R��U�����]L˗|���h,��¨�g�-��{7FQӚJ��7�[hW�� ��,g3}t�1M�U.��q�����j�H�^aw�|§�
E�:4nZ&ޗ����n1�:�YU�?�j ��u�OJ����hdS��,>j'iYg���J�9��ʹL�-���{�F�dDn����A'Ѭ��\`��q���髝�胉ϗ�Ǣ^��å���D P���.�$v����K'F֦

*��(����x�Q���W�놇<���H�N*)��<Z�X��rvE��S�����H�?���RX$Qbk�q�р���7�6��(�a!��«�(�Y0F?�6Ve������T����T�_������c+ �><�@<�O�[�{�t �+T�#��$6m�TV�s��Z���H�ӯ�8�����Y�3'��D\b�Jb����{�a0u�������Ѐ���L=�|�L��5~�&�X���HЮ�� @^]^�^7��6Ra��:^�1[{���^�ǘ/�Z`�����&��8�9��a<�q��<#�A �M%��� ��u
 QD0�dȁ��ЁK?�5�?y7����z���F�HL���oe���*��r}|�(a��<�غ���ъ�1��O���ծ���I�m=��
=J|A_W�6/[YE��B�(K��1�ɵUg��Y�(��G>��J}0�.
���!t��f"�����PFc��#c��ð�-R��=t�f O��$�)+9Ԩ���6��ʄ����-��\�\ Q� ���"ghjj���G����~ 1b���?���s��'=	
���9x�fw՛�T�P�>�c��3 ���?�S�o����!%ٞW�W6�B�>��)�����Q�lx�Z�ic�	�Q�Iu��_�5���z��`�?���:��x1	鶕�vQo�N�S��� ������H���D�{�Ms�Ї�6�� �s�Q�����^��H���i8�K1��L�+���p�Y��?K���R�����7@�~��.��͘�)ȠL��4���N��G�o�hI9���15�?�<l��0��"��W�M���N�[��7��j#l~�,�AfKtٙ��Ȧ��}�>�3��7��w(�Τ�_Ӽ�˾ye�Z*�hf�W����t��X@����_ρ��Bar[2����F�u�^��f0�b�^�K�@9aY�O��z���v�
��5�G��m�7���H�ޑ�Ng�$���Q����6���N�|,4�9�y�)����g�@!=� �a�ja]�u"��Q���L}_�2����F�L�Ѻk��J*�M��8O�F�����jW�YG�E��¥�)m1¢�!':QA]�okŹm���fC/���_5��� ��f@�n��T�ɢ�u"�@���b='W?����Qwx�Ȥ3j$αͧ��YGqV�\]7���L���1�]�):�t��).�����f��u��Q�D�*M�2��.��eg����F����z��'v�ߚH_�Ȍq4��VF8v��k?يzYy��4m��򝝪�����aC��+�\��O�����v����&P�o�2�ྫྷ�3���j�����1�'��O	��a�lq�{��sfC���ݾ��sl?`�[��(~t�<�Dm<W��ܑ�u���"�OS�����O�f�n����Cn*��z�í��nWI~�;?��<�e�!Иa~:@�-8��[�;ڶU�]�%E� ώPJi�ZJ?�Gq�,:^���l[Kj���W�d����Z�so���A���������fG�t	b?��w�CV$6�J��^_^�H�qmG�ܟ�v4G~�6��{9S�&�{z�]���u�L\��y�׸w��!�ò�[R�gurjr�=��(��mYYs�0�z:U%#(�t����pC��s���"�P^�n�i��<-Z����Ax�s��-β\����&�v�T����P6X��"����忢��|Q{�4h�ɂpº�ֳ\�@�8E�%�ZN7���iE�LG!��H.����,�x=ǴUO+E(p��Z��<ո����F��7�ₐ�������	5{�<UEXs^-Zrf�p���� ᘬ#.�!�Y�����2�=V���y_Y�=/������T{0���P��P�#R)�@?�=2�>6�-�Z�Z�d�4�Ԩ H��V`<�I m�3�#1�:K�-3x0��.��	XWd��[� ���n���S�a�I�;���E�d��7�؎��Ju����ٚ��NM� .���.4ރ:�h���e,ҧЯ:8�rgڱ�Xu%�-M`hr}�#���x��n����,\O�-�LIb�����
�n��)�G�#���0D':E�F��V���B[��}�T�oLA���8�����Z��IOnz���j���i�o,
����
�L������0��=�_Zۙ|t���BN.<�,$�_$�0[��j���ܢ��������CY�
uj�b�+	-v��������n�ފ�ms½�s}�������˞�����5�9��R%���t��ʤm����`���3��4
�Ԓ��S�K�	�zl���E�đ�V�X�A��eiz6d"DMg���<q6��M�"���Zq���l]�,�nBA�m7��(P�������E�gNp����M$tHSc��sY�!�7�Y���SU���1т?߬B�^ Є��k�ѿ��C6QߺBFf�Z�J��0���%4i��
��>��IES"��?���|\jo73G����1m��r�D���$�tĦs���r�"����3�-�>�s6��)+�T5I��
j��Læ"�~��f^:Q�K����͗pԫ]��H��u�r�ۺjJѶ��.�k���:�C��dI7�Y�t�FbUK�C�3�胃���@� @P�W�8����\��x��]����d��a��`xL�nfWU@�x�6����Q�:h��͜��h[�W#)��x\Qj�]<���4��(I2�8��)F�0�2������FĿ5L �-�8���J�lv@��Ϥ�"�����~���"��&�Q@���Q�����W?�@ ���t��IMb=�>NQZ5����gB�p<�!X~�1��s� ��%�,A����<-.���\-��_U�����@1�dU��JY��`���sX�};-�m�S���K��۾W�B�~Srũ����U���FG1���������3$���Wc ���Z�N��3ɳe�=|b3�޲{q~�|*�ҳ�*l�:����\�H����ђu��a�F��&8�t�S� �IS�`�Fn�n\'Ga�g�,�9�؊	3������k����RX�3�������O�j���:�粠���4 �m)���`kH�J4�����g H��)FG��%��|7�zl؜V\n���G(��'y���N���2�S�5�����^�A�4R���Z4�F��ߏ�ʞ��~b�z ��)��s���-�f�4c�_Ewq;��o�5䡦�}����D�q�U�@��(xx�=Y'1����bTB{[�p�LQ��W�8_��Vx:Lՙ�ڥl����%�@L�膷�!B��ȕ�t�!Ƿ�o�)��p˛�;ֳ̕�25~h;rh���%�h���(���Y�7�)�1:�N��ٳ���F�u��Oؤ�7��%��̊�%�9A��Y*����3ɖ��,;��x��Pm>�u��РxYU=�kF��NۄÎǱL�x�HS�-s�C�e���|�s֪6�xe�1'N(Z�!"
�Ҷt��:�8DwE'�舆!p�.�˜pTq��>h��X�\$�"4�1��˿�,��E����Ud�>��}i0�~w-`5r�e�an%�)��;�D���OK>�e&/�q������x��11	0퉊��tP�Đ�%訠��l��];oBE4&�c傲:)
��F:җڭ)�ר���Ti���o@B���1�(�S/�)<�0���P*J���g��W�n-f�"C}���j`��$��"8<�|��?�pNsy!:�HW����:-�1祐�'���W�ؑ�Ic�U6jr�`��p!���^R(�G>���_��a����f��B'����K?VK�oy�a��ݴ
�B ��B����q�y�~=���} �,֛�rY�2O"(��Fo�Z��-���b΀}��\޲"�y_$�7�"[�M�T�=������D>zL��r��ꔡG�M���������'B����1��.R*9mf��^ 6�v�8��e���] � +�P���Y�v�Ş�m�ДX��������ؽ�`5�_=^���~��z��<��w��LhFpa���ӭ#�PWF���W���q����7�-�g���)f������ ���#I��7�-����� YG���E���8�R˚j�����,e���(�B��im>a�dM�`IʚX4	<*v]5L�%b\>67$l�<�N��ovJ��՝�R{O+�2lM���83���6e/���{O�>����d�c�9��E�FF�m���i��#������:��`��:������Ѽ����3���8��|�,`d����:�\"eˠ��M��Q�]���S
�!<�	Be&�[�2?���Т�̍Ö��b*F�#��x(8)
���}D���:Y���9��.����6-nZ��f9��s��IV�'��z+�t�i~i��By���G|�����l� ������#PI2�p�}V�q��C���K��(��(�W�֝�N�-�E��e���l����'"EM�$ީ:f�q�)�����B���s���	���ʹ��B/u�Wt��˗�6f�;�֔RGkW�����0��b��W�$;�a��b���/E�Eϰ5v~ʼ������jB/]�}?ut�l7J� ��9FV�zD\���ҭD�'��j:t�
��`�%�����a ]\	m�oG5>2��:=�Q-W�s��`��Me�2���%7�g2����ƿ9KC.�e����� {ڵ���!v)0��w�0���:���a#�q�I�Cт�n����7!�����^�w�^��$g�3f@����[��u�Kb����)ъ
����^'����mpX��7�Iqy_A����)�HnoN*&n�'@��sB� �1E=Ǧ��-���g!*>�3���7�6R�B����*
��-�ۆ�����2�!���% i��вZ�1(0�R�]FA�	��^wRU���k��ܛ�M����-ќ3q�*���`ܰw6����Kԫ���,�W}��ϕVU~<�ԇ��ϲ��y����v���W���rI�N���P^��_�Q7����71��Ll�zh�פ�J�OqR{I�3S�P��}�5�b�����/��各}�Ѓ,���{Ɏ{��~�I:��B=g<�[�^f&S���PVn�����D��=���x�%ⴠ�΁\Y捳�$:�)2z��z1>����k�������U�~�gv�u���M:�Qe|��D��� bC��Z 0guR]��'NF�˙V���	��Z��(� �n�y0+Q�����o���XD��̹,(җ���D1%�*А�9���[ӝ�B�i��h����$���Y�(����+�>G�)�=��3���3�ipg�L��
�X���]ُ��D�;+> E�1^�@1������_м�������3��F��yA�Q�[C3=.$��1o�x�y
��'v�q06ҭ��&��/�p�$:2w���h��e�I��A�ظ�.���<w(X�.�B�F�P;(K/�z�6��ӄ��HG#̗KW�{2�H�,����{��
(%&0��7�v�D�-��S���0|ʍ��5�af���߁W��BhDcUV���:�]	8�I��=��z��0]��'o>����4�7�Bf��Y#��I�E��oG�5�ˮ]Z��:��wu���9��Q]�����U��r�OҪj�3<Ty50ԇw!����$����OK'��	����NC�ٍ3D�+�`�9ˠ�1�9��9�;��7����J�Sm9i>,����V	s�n��h���3� *��u[��ړ�i5	W�Ȟi�C�E�=�ίY�)���}��ZK*�֞G]_��|�&�v�G���X>ڕ�*��g�U�J���w�X;�)a`�X�i
|�{�i��3[����|�����`�sn�J�9� %o�U��h����f@dпU�%:�:�!�#0j�Ҭ?r��Uo���2�Z�"K�eN�5_�W��H�AI*�+T7,�z��� ˩vWr�J�E.A�`���yi�=KH֍��S��G�W:�����]h���:�x�/��T �����ܗ�b����
���b	�M��c:�S6�}�|F��#��FWc#���W��=����$ׅ|.D1�~�v�XdP���'xI���!�0-ј8�4 }<�=�����8���N�){���2<`�+��fb�(&���1�h�X��u萇��9t�Z_��+o�3ur*+��w����\ �����
��D/n�m�i�B�܂=�:�׻KV�3\�F^�:����Y[�K��c��;-w1���udh-*Od$�dp#c3~ �:~G�MJj�B�e�(��+c��[�ނ��WW�D|e.~��g�Y��)%���hۨ�W�~�0���gI�{"R��y "�M'���u��;�I�G4P��q(�;�vV��B	֣�f;1p�qpO������i�k86����X���L�&��[��/[�����q~��0��:W� )e�Kvw�0;�,FR�8��
�D;dۅ���Pp�Z}�9T#[Zl���K��5���Æ�:%v�ݕT��j�7]u��{7]t8����Y��)�V^��H�%qn#�Ӫ�+����^WS�G�c���)��Z%6�,�*��T�IE��`��$7Hw��-�o�t����%�1[���3����@}S��HS��?;�(;�+|u��5��$_\�! �V��D�h�?�{���oi�)�v��5���@�����uf8�D�/� NR����<�~��ץ�������T�,�2�J=�>�<��I\�AϢ�S�0���j�<�w����K�A��ӕ���ф���DDe�۩���e&�k�&2�I?]��|o�{M��t��2F�ͤĉ2�� x����m������xE�Z�������ر��t�
��@K�0�!�GXk��G��L�LE)A�� k�Z�M3�/�}����Ul�%H�+`��_Y�LՃy��ۡ�J8ˠ�ļ-���ƌ��$���5�՚n�GI�g�<X�,�Lrʸ�6&�X�X����?Ia��(�_� �ު�Z,��������W^ �##c�u��[��W\����*�Ie1`u�L�5@g����L��<β�-w2��0%p�oϷ�DiKYY����߾����a��)k��T\a\R�5�	�F�I����a���!�H�~��㏘=����0����a��)DQ1������~_�3p��^˯^��G����DJe�R��g~=���֊>�	�C&�y;a�}Y)~\wf[����J@�%�������o����\��JZ�u����Q�&g�*I3BFW����\m2_�n�XJ/��R�������}F-����������l�p�r"�����-��[�8���³���:j4�c�`٣���,��Ms�7"xgH^��nM^O.}UM��WPpLu�F+i���h%]��̶8�%���l�oNV\��(�yaf+�.��a�!���r�)�,8*��� 2�SF���ޛǺ�Yx����R�_+$��J	h8�۔	�s���m$��Z(�9%ӊg�
~��=�T?C���qqL�
(8�-krph峓�8.��ye�UBj�n���G�Ͽ7[�9��ڨ*fޟdk
�ޱ�����E�:W����	��J�@R���V�ˇ�8EKI���&��*�؅W��opz}vϾM[����:�R�'$���~��C�&fV�Eډ�hs���Ô���U�~�%�p�h��O��i�@��-UL������B��{'�Q���ݩZ?��8C�
�����:�!-g�uf+�!���\L:��_p"g�m�<)���<��ݾ�ܯ$b�yO��!?iK?�=ZH5z�N����Yw�50[����=v��˷��o�md��l�]��~an��{�/�t-��h��M�J�7���z9�wC��Tuw��U���YEiv~
�X̬���.^��Y�e��W<�[��aS`�����x�To�5�:>l^���ŷ?��c@��a.���!�H4&�@��ai
�";ƦYj�:����%�1����]9*����u�>-�� ��<�|%yؾ���Bj��M2͎�Se��r�ܻ��z�+�2?ٲ��I��v��j�!��5Zu�g.Y�
 ���3x���΁dS\NU��K�N+9:���%�
�:��fm����آnMK�R��j���PfP��^��0ؒ��vj{�ő,g4�SQ���b)��(؝������-���Zc�n�{��?����H���<��8u�Hu.'V���d�P;,H���foV;"$P�hxңpN�c[�ʂ�fldc��,m@?mn�ְ��vBJ�oq��|(��u�����=h���*�PҶ�Xa�G�5X�9�d��b�3]F�H��/�A�v����h�S�v�G�����ᝎ-"�L=� {��S�Y�ڌu;�۞�QG0���I�M�&��6�"�)�ۿdŒ�V%Y�9n��Q��|�+�5v��.�I�V��2���^6h�� �l��i*�~`���H�I�ܷ5�vwN�^�%u��wz:u��s�ʻΩQ��oH����R�{�������ɑXA�b���z� ������op�C6��3�ܻ����O�2���� �\v;a�p+�U
ۍ���HM&�|��&~C�+�PVk���[;o���L)�T31'��R*���'�冾㗾x E���b�K��=N7���Z��c�ve|Fq�?�b������Q���X�Z�����~ݱu��e34�<?��E��
qq�t�"�t�Qn�WR�{ܙS�3��hʇ29>���X&�����;�V���Ufrg�D�7�����a�V-}�'E����BV߸ti�9z��w�#W��am:���E��8`���)�qY���ɯ���Z�n���o���R���J�l,�OI��	Y������phL��7,���-&�ʤ�m�lT�ki���<����\Hm������<�U���\��|�K�{��ZY�Ր}�2y��Rme ��S"\�V�~�дN%����	�QyB`�B�ֶ���	�V����x8��\��v-v��ԐA�V������$.D�����M�׿cl�(G!�.{.}�BX����A�p�d�uN�ly	�sB:�N��P!��:|"��Нfi���cL�Y+���*\U�P��1�]S�a���ɉ�HGX�j�9!j���p��KQU����T�ۤ=��=A�ޗkiJ���D�Q�<3&���y��FqW�k���G?ŏ-V�Miʦ������O�6V�c���*�$I�o�YW
"[��~±Phu�G�Li\ �W�-:��팰fydTb�y��1�� �[UM(l?�p�U�	]�@!�ڴ~��6,����p�ingR����h��8'��	�Fy�u�د�x"`�7I��V�  {�b�� �N%a[���+J-=�q�4Z��}D���0�fy콎�"_Ӎ*
�x���	���1Ӽ�_�A�\�p�;��٥mg ��ɒ�{�O��Vh��&%��J@2������^s�w���{�\��;����V)��f���]�-��ۊ���1f2�X�����f�7͏��e*�!Ń"6r���A���>w�~G��Csy����
����8I);|V�k�Dkw"f����YA�2���OX���6�M�S{<��R��-3��bD��[�}��� Rb�J��Ҡ'����lh������]��99�/S�0������ԘAf��T���5c�h.�͇bPq���f����_��P�='6����|�;�S+��{[ˍ95�?��S����� �o�g$�����@>��v��Ȑ&���)�MØڜF�vC&FB,�w�3X-qK����}�P��԰�h�q ���Z.V���B����hs,�7�:[�-�GR6;*�>ᾕt�ғ��^�!@4RJ�P�@��H�L�L�$���Nޠ�u���g�;�ˆ��̸�&� ���O;5*!�,iտ@�I�R+�����u���;!�*(α�\����щ0�B��Kq�"�zv�9�>��Z;h�q�p��Y�h�P�~䬏ߝ�ծ��E��,6�rL�S��^���f�6LZ��0$v�����:�v+�Pd�.�h2�?�_X��,_�L�r����z'��6w�pgtս�Ɓi_���8�,ʭ`c<�8�={�@�-�k�F�,5w6"Ng���.�Ƨ֟�?UX!n��:h��'���K��9N�y�����#`��$P�/�˶L̐�t���2	���r2�ʿ���q�i}��upK��|�$�-I��"N�ج��1E�ܝ\��͵��*Z��@�,C>Q���S�u0�2��z��k�*�5�mԟ I��*s�S<�Ϛ���A3g��(t*�Gg�VSo8�B����{�e@��|f���fI��� j`&�����'��Sie��
=�w�P���o}��P�νa�n߶��7��E�;�MM�̾��(���`0n1��}eu�Du��X��Պ�i�c䓥�*X�N���Z�4О���2���а=}q��p���*Y|PYn^�����������?���D4p�.��Y�ຝ�œw�� 5A*�E�����Z�#����z��������;��fm�c���
��ל�o�7�W��"]_οc�*z[����4�������HgJt\�[+�(�����<��02ٯ^^2�:�������à���J?������R���a��"����+G)>�.T�ܖ��s�w�$�@b)�{�"(�\>�C�}�)����@oy�S;
~��6)_����͐�,�U��@�̥J�(�}�é��cTUL�o'f�&�I����&ͫ��A�Af�K���İ�5C_�/�9�¬���)�;&������`X�S��j���%�sg'4g*������z�^���d���; }1r��2��؃f�bZM�H\��.O�9����X�[�3���g&׻dL���P#+(A�݄�OBD�V�j�i0��H{#;�`��Q��1U��������a��Nn�`��r��B�Uܡ�kU#V�VOn��7�K�]�p}�2+���[�m�AO�,%Ҧ��
��>`\Z�jK^�`�e���\�M����	+�h��y��9��
��lim��>yc�����La6��3E�='5���v��e��d�7���U*���N�p��C���QK7i��Y��ޣ=R�Hӫ#}J��Q�@p�N\!�L0���-)�ݧ#Gۧ�U�A}r��V�%�����7A��v-�� Y�X!겁6'��i;Ø<�ONO����3�YN�Oߙ��X�bA4+��5��̴E�� �Va�g�@���ߚ�$F�y	��a���vo��i>y����W39����n��c��8@Wl���;=<����_��.����F[Fu9͓����!�?k���.�b��y,T�Ju��C���<@	ns��@�{������P��q��A�,1O9����4l�	1�ʃ�\�)6l�$�M�	;͢��'̂��mp۽j��:�گ  ◞��v����J�tgt������7@���O�|]�b�HJ:����25��ݬ-�4T�F���]�X�w�pFh!�Z\�*5�̞���a!�hO�W���^�	Z��e֦����Y��V&7N�)��G,�}��`�G����!�-B��\Pzb�\<�F������h���@���Q?��t���B?RѭX��r�iS\�O֞ú孰@�uk�P��X����>Vr���C�d�b�G,ѻ׿04�&r�wxUº��b��j���߸�UoP�_�i��J�����n�K�����`��jA]'��ٺh�P�ʺth����u�^f�:�4�!�p�19���Ȩx� �������ϲ30��)D�I2�ru�P����Q'�(��æUvU#$�����>C���*;�n�NOj/�̾��͇��(����d힫�S,j0?�}2�P�ߊ�pBV��ϩ0���}�χܔ�{f��W(��H3/(� �+�����z�*�H��R�GT��eS��4�Ha!:(�ym�z���n+�:[���.�ջ����h��Q�M����/��J�Z*^p;��.�4�����~y��d�H�g=Qǫ�E\���*O��v�fI������Ҝ7ɳ�mB��mC½�ǐ�%�~tpя�'���#�Ƥ`F�$Ձ��d�Ŝ>Y���
�k.�˳dK�Юq�lYG	���
ă��U��j��(�|����/�	%K�jy����2���f�kO�+��߂F����A�����p}����N���ۨ�<jk�]�,���]�d�G|+�A�Y ��d�C\����L��A�GUW9�Ջ�e�H�MT����н�A�`"�v�"��؆E��pM O��6լ?���r�!�ϯXأ�d��bW1li,����=C�vW�h[���mc��a�qoB���5!���g��J�n2����:���kD�L6�zM�@����S��*~{`yX7�.H[	U%_���|���r	��dm�":��<İi���3�/�/�_?�ڐ��a�-�&CM���!7ߥc�``*܄6�C���d�.%�Z떗f�S2��� ;���x�3S�_�"�R2�	���D
�9�]�����+�� ��j=�nX��sn��	��!0��ѵԌ�z�"F`�����ǇM5�Ή�9�V���#�׾��@���w�5�`��m4����J�������ʅn)E��	�R>�bp0�@q��S>��O�J?�7�L_N��t/P�h�U����ᗙ]�^dXa��ߩ_F��	�cn�6��S��Z�J�U���S�Y���-���WK�2�L����|�ΔBw7*�Jʐ��/�e�&�WR�鏙ydʬ	vۢ|V
fb)�~~�\=�G�̜�_�́{�ϕ,�~��-4۔۽����Y�����NE�l�&���T��Tn�۶5��&
�<b��*��l��l_�#mƓ!qݖ��H��#�ԑ���k���I��2p��k#B|:�V����K�L����Oֻ�*�`�U!��f�M�D�ﷳ�X4�F���0v��s�y��v�i>fLʪ�b�֖��;ץ���~:�-��x;8�
����$�n#�N�ԑvĊ�;FZMC�wx�m��ǋ���@�e����i	;X�Gظ�I�&~��	�9/&z��T�)sO����Zﺦw���B'���&��?�!QO�rd�3��w�.�ޔ�T1��M�ѭ)�k�4X#D�?�w,�[Gh��ԉ�aHF�@v��>@@J��R��!h��)��Q=�������ç���(��
Gۼ���0��8HA"�k��=��j���4���	S��i��50fFO��ou�m�a�8^D)Ob�I�����O�*�u5 ��b'��W����뉙zG<����L�2ʷ���Y��{��qe�ce"��'�$6-E�p V�P{���&-�0�����b�N�&���<�5��e�`������R�wv����Y:�/g\K�]���gQ�&-������ �25��i��'80��q����>��]]��H�6@�Ήj0�Zt	�4���"u~vC�>��8�?N򧑹o�ޙ[$�����k��Y�-���F���k�@%�g�Ɗ���?UVr?��/��G����n��#`��,�[o4��Y�. ?p�����"�����㛶�����I_\m����[�J��w��@*�W��Ċ��n�酤sƸ�k�V(^ ��oh��E'I��ĵ��a4�M�k���[�$Nٮ�}�u܂�뿭��?ܪ�p�'�:���P��G-[eT����h����x�HךYP#E��c��#(�-��W��w`^�˽�H�}U#~�h/��&�,��a���D�n�Y_:� }B]#{} lV��Í�Y􋵒{����p^�@�=��e�����6P�_�:����J {	��p�<�;��ܑ�?��U9��wqD��UX�H�T��TuCa�f�.���|!Њ��a�2��A�B���G ��Ͱ������^N�g1'm��VFY��.fPAʠ���u��d%��\>뿌��W�|u*pd�EIT�}E�ڷ�'j������ $X���l|�s1~�SO	+�.�k���j�4�}���/R@��A��w�s͵�}��Lik��'Hy�`�F o�,?���پ��>d�Ñe�׀0ǋ���y}'�^�2�c�چ�z�o(��{����yqg?����zP�Z�
f�4�O���ק������a)0����HEl�|�6�jz(�'1o�+9{��pAE[�����n��2�C�E	�i{���Ȧ���q�mI��ѹ�hn���31
�ŁYlN�z���Y���H��7-�=(�v��{	������|�9�6zFje�w`��@ߵ��Ro���^�n�>ki�!z☊d�i��B�lD�45�l�Csuh���,OD�����<�g�w/��Q.�l�Q�
s�x��+V�	���t�{kb_�1�l����?���.D;0#�o�7�Ȱ|f�Nf'B?<6M[��r����ON�V�f�f��R�l�7�'4.SL�n�Su�w�1����qL��{�tI?}����N}�1���Q`2ܚP�)��%�B���{��Ա��k�J	0Ltl���q�Յ�RH@4�́��FE�Mu)`Z8�G%z8���sS�̕��[�T�{n��C=��bM�Sh��CG��(Qc��d�u�o�g�b�W3w�)"�#��1�b$�j�b�3F����E6���e<y��R�)b/u����}�,�*�X_?����HYԞ�pO�퀜�.\�I�ܽta�ٕ|ɝ�<�Ȝ�=YlbĀ u\碹\W(�x��F����~���#�V���C�઼�SC��,�e5zS�%�l6#0J����� �n�6%��=�<Q�j�aW��Eg{R��<eΜu��q�e5A�
�&�EJ�ƴ3�צ����<-E��@�<z����U�H��,mQ�>�ǢBX�l.A_w9�/��4 )ݘ��w'����ޑ^]K� m~Iz,�/[��8d��xca�f'�τ��3�o���=e$o(�hH�x�%t���*@�	��F�#���/�B_@!����ة�蛪��g��0m�����hɏ�|߹d�(�`�,���к��,�n�:g��<6hWXb�Y͝@�^ .kErC)n�\.'B�|kL���`O�;0�4��Q9�C(�b
���!3Ch�(���ĕ�`Ag'��5�\=�KZ�� �h�ɰK��Yy�G�LZ�np6R�y�e]��D~��&��L�b_R�Ws:	5p��	�f蟉��Mχ��Ę�S�0������S�og�qJtVr3�D���^���t9+|TOQ<���b����.,(����X�6��[�`��Y\��UxUL�=N����ʁ�/~� ��F�0a�\Jƀm�A�������=�i�mN����-���*�fYURs�[⮆�T�F?��1�
 �c.ED6� *�(���ۼ.�sfD��֐DN��XP��އc<&]��;J$4x���9��rr�Na�Y��ݝ%>s�9��p��T���&���qk��K���kG�dR
<�`* '<���E?Z���^���K�&�(���LAػ9�QLn;��$G��/�:�a��v���f����[J�xx�28\xMYנ��d�*��\����S���#�4��3�ݡ��[
aQO%�>�� �B��{<Z�!�[�!!	4O� M�Hſj���}��.C�����Z{/��NdY+�k|���)G��G� �����0��C�2�Z%О���1rJ���'��	�&��\��0�mr�T���{��P�S^����R/oM%JO��u+��V�t�9�����"�m�v���V�#�n씔��2�����hA�Q�`�'�J�Z͇fm�%�Ea���	6٨���)-��tz^�P��1wo��-���b�&u��:���&x�ׁ73OfQ)�#χ���p�ٖ��		#J�\��~�I9���q� ��M�\��'�
"��Wٺ�����TÚ�����n�tT��Ol_��� ����4?Ti�#��\�g�'�	���;$~S>H��H���)�H�g��4B�1��^�c��M#������o׏����Dj2�%��-�.�o��+��m��u(U2�-|�����6*%SM��g���h��F�mI���Ym���q�Ћ�%J���$�W5�ݮ](��KFPjC�eѩ���؁�y5���+U'�>�%]�5��ֶrB_��%.�Ԑo>p��M��1 �k���b���aR�3�>E���7�^�����?��K���|�S����Q=���ߑ�O��Z��Ri$X��{{X�kC��]R"l���X�W�5<�|�n�H{ZY��I�|�?y����
�q����m�f{���P�����I"������_�5a����K
\�p~R`cvp�a���܀���h$M �3�A��og��\\���.��J�����x�p�� ��nG���s�ݥ}����Hb"�y���jX�����U}�c�[ݻ�KV�����:�6��#_�$ԩ���r���!;���2��k�+�*9X�$?���(Z�o��)�h�<��0�=�ӚKĭhC�������g��?�iē�,���W����9=��o'q��E��](��N���K�� ��j�^=b2룎��m	vNp�}+��h��|vi�DV��R,2.�K+�t<]�W����WR]p7?��5�R�����:I�e�x���*���M¨��A��œ>����Ǖ!�����c �	��
2ڒ�#���A���"W�hzH�� {~͉�
����/v��k���ٌ�\�DeoėE����P[�s�v����eqz
��bU�:��&�V��G�������� 1�*��>�j�w�r��C�.��3M��t	��w1�#1o�>攸�I9�k�7����.5�h�>���|������(��}�ɳC�)�"_���O.t��~G�\Y�m�4~�D �I�9��9����G�b��h��OdV�� �,��粪��䀆O�6+�\a0A_����_���*�Ro��؁<�{� b#0�bH>�PKl�m�߂&��I��A��ipǰ~4`~��P�6��>� �C��ȓ�	0Ȝ�	�,�c��8/�qAG4�n�H�cO_�`].Lb����&�TIN��O"�n��}����N6U�����5=�:�HIq^O��|�����)���UDJ��^��K����?uǫ�0U;�cm@���[hJ�o.��\P|)i|v�����He��a�d�
'�^3NF���g�l��اL~s��}N��.gB��R���
+��G�2��,h�����85k���wuƊ#j_�~&����'�ĥy`�lLju�!��ʨ�/_���O@2x�o҆!mr����J�������Zi�Ʃ<4v6�k����'B2Fy:e�7�m/����+/"J���r��~�����j�Ftb%<�ԧ�D6Ǒ�S�ކ��aN18��a#Y�;�A��n��%N�F����m̫���µ��߆[|���I*4���E-GLy ��kg£�%^�oX{e��G[��������@~$�,4�A!���{ qrR����
zͣ���mo`g�P o%P�2��P��Oi���'m!+���/������#_x6:%�S����R!>{���q��v���{޺�Y_���6<	H���#N@�����2����=�+�H�߷�Z��z�����IG��-Ū/��$z!���v9\���l��Z�у ��W\��A�$oK�(�r�8K'L��#b��	�ܳ/d3�n�^A���T\K�.2�޹'\AWYF䞶��{�{7��!�8�v%뼿"����%	R�"����o�ҽ�o��j�Q��#A�0�}��'�a�}��&[��)[� ����_խ���g�~>�!?Nw���R-��%`UU?e�C������@�8ٺzW���7��ƇeJ�_�r�	�Ґm\��2Y��'��^Pk#T�V(T����&��V�8�A��^Hj�9\+��ה��X�Ғ��Q�I���"�^��&�R-w�N̘�&ݝ.s"�|�U�����~�<V��{����&?�^���\�� ���89�݆����NZO&�~vO��	ʇ5\��W��<���G��TW�H��_���[���~��g	��|ySB� }+�~��0|�H$j�OC	��jp�p�UXP�D� �J~F��^W2ׇZ���� �\wj�3Y���U��q^��k�L����uŢ�_�v}��R���'=�.�޻�!�T5���¥$��Iur���F�	����vѱ���@�d�l.��-��T�.�/�L�ɩ��0��*�#���$qK�ʙu��ܠ5H�0��\����kRt1�$U�1u#0�"f�]�/c�?���cZ ������x�6�a鹗�����O%.?��5'��#\9��Y
i����ve��Y�w������l��'Y�AO�m�E�\��ij׈��R�ʒ�4�n�PYܖ��O�.뿭�C��$�
4���π��he�� !Ga�������FP�MΙ=�W?Q���Z!Ǳپ�Og�[�CB頑�C�x�^�ҝ���LJ�����R��0L\�
��hB�>��9t>t�����3.��j΢�,�^c#�Q�f��r���Bd	8n�(��"���7m�U]�&#�HzEl_~ټ�4`�8��)(�0C�3�������D�����D�ai�vx�Q	P\ᴗ���tm����B��E�C���C'�M���U#p�֖�y��VյS��44���X-�H5�z��Ҙ���pc�&`8_��^����
���z����U���3s���Z��;\�\w��VX=Ť����⌹�Tc&1���ux��Q,���f]�FLq��7ېG�<X�]W�L�����t�$RJ��i:�����䟷�T"����pa8������5��:�_	��6�o�L�S5����=�B�/�����P]� ESze�'ӠCF��\"�(�k�yV�{f����I���L�%����TJYt4�_q�\o)�d�KDq�qH�.*��0�#�L��u@������������'-��Omw��
�v{�G��&A�"��ϊ���)