��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_Kq�n��XaR���(T�,/=�1Jny�/[*�����Z�q�	cǩ~���nv�FmC����[��15/F�?��.���}��"d�D���+��O+����d�HZ]�I_F��4q��w�5����&�NJn��K�
����n<���&Di]��vy�]�<U��ո�|sLCK�ã(��9�S�E�<&��Eɋ�H6/���>�a3I_+X�A$�q{�V���������n'˜B>���X��Z��>���&c왛e�4{`�kJސŶ�0y�{�}�O�혝�`^Ȩr	~�@�ٙ�؋��� �uvux`��@Q�=������>=�����]�{�+����R�3����~#$?��l�Ę�aɣ�lO�s�� &�O�E�7>����RL�<�|Ӵ@ҔU��S��|[}�:3ג*\��-0k�^Jo|�������'z�[�v�[���JJ�C�΄0@��U�`���U}TZԄ���9�y��
�A7��e�fCB�U^j]s��uݬ3�08�������լ��uU;�m@N��\d2��IE����ۍq�ȼ��_HP���	R�aײ-�/�-Ź_����v$ Plے5�7�f���Nf`�B˾���N{e��f�(��[c�p�-+v:OQ?��ol�At�q  ��Y�.��[2K�I��ܙ�,h?�0fNZ�~���T���|C�O��QV����\����,k����- ��.��4)iTG獩ɿy�O�1�<ª,�alژr��y�-��'����?�JD���( g�^V�̨�Jp�%] ��#tEo5�	0����5�����%�p�>5#*|4��;����Y����.�7M}(&