
module syn_threshold (
	source);	

	output	[15:0]	source;
endmodule
