��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�YM�C����ion�W# �V�Li=��?>�2Z=p�xP��� c�5}� ���3�}��j�o����^�ࠄ������G���P�z���7R�1��I,`�Bv������d0&���`�\3K�j5n����+���AM]��YV�=|�ޟ1�8����v�_Bc&�F0�\�q[�b�H���~�4-���������ΑQ������|�
H�X��������q�aj���Er�T7������ڝR����� ���U���,����U(�ʧU��'b��r��εoLYڷ΅�H��p��A�R�RF��Ҋ1:&��Yuc|�o�oQfTo��=��GZ=�-�j2X���֋�Ƿ�N1$q�9��?`�v�HW�B��8��p���)4Ǡ�Z"S��(��}�S�%�	�om����e�3�{�Ͱ��g�V���eH��$��#�����6O!/�4�y���]K<(��ZI*�U��D�����ȣ���2�23l��0i6LQ)	G����!B�<�8�v�*8 $;�ұ$:{��t�B:��ǣ�|�VR�H(X����n�P�P� cU#i=�>]� ��H����� 0����ehݞ'�A45������\:93l�*g����-y�W68͵>��Pcu%�0`7u�I�S�!�S����}_�'䦢�rD{��^p��<N/��.#z��R���	����c�ɥA�Oj�Y�˸�m��K���ٿ��◛r{j�#*5͙@��%��p�jF�p������Z)�d֗W�k����jŰJI��������"�V�hG�	/��q-tB֌���dOy���ۻ�����>�(�T�����I/�,|�	4��a2�\\���Ht��>v��"��L�6����Y7�����RD��1�5��%�$���gjW�W�bO��3I���q؇��&|�������@'�～k�k�QY#
1�ĞzK<�m��n㸰����ߖ�i׉�PQ�h�˂#;�X�>ɬ��$U�~%��()����؟mL�;�	g�aI>�e]� ._�}�hh�9U�UN�)�Nr6��5�b$;�<��ߨV����47�!��z��5+]Kc>]x�E�l7�!�|wL4x��/9~��UI��&�-���e2X˙��l����O��4�sL{pz<W̖��С��,�|Og�l(�aj�����)(}.ɝ�R#��u���agK	4�7���e)3m9O*k�jr�D�����D�1��ZS�Z}/
~�0Dk�<�Y���E����1_
־��R��L[��f�6��ϣC�Rh&0������YRm�p�R�~IBT�*�P����fߝ�n��8�6�\3ʺ�v�%�6����ԳM�ޟ��3���� 0��@@��I�\R��#!�moᳱul��"b��R�5���ڝ;�K�%�Wr��}
��t͒E9��rtźv@w7,�Q�}��6��{�6Q�
�L1D$�ۜ��.�K��59��7t� ɣ���2X�#�û<�8������g�������j��<
u��>�#`�3��#P�3P�O�%�e�X��V%�U!��F� �	̸��ь�cs'�;����x�=��� q�������˫�㸄M,6�c��׽�� �S��,�GWps�
Ĵ�*P|K���U�V���=��4�^�Y�ʛ܊�N�����)w���.�У٦+UW�)r�5��i���c�{h�Ӌd//��r�A�m"&�t����[��0����σ+p��M�Ƌ�`�>"��M����������_���)�g:��h�D<@�+�X�| �Ӆ�%�HM=rN�$���c�@�gf�f�e�, �9�з��G���_�6v����C��a��6��Z�H�6��p`I	0�2C��_^s�T�.=������F�z�^d����-B�{�6~�-� �^���|��n�"$����L�q�`x�r"��Lq�c685��W��|^��� ^Ʊn�(ȤC�N�Ӝ&��:�9_@�-�7����[��p��e�9��z��(u�aM'DT��/�X6�H���\0�}Y�����g�έK�*��c��u�Q�ˍKi5�ȡ��#$��O�.��V!�
u���Tx�>�{��u��(�"�Oݾiy���%�;�?cc�o������uN��Y��Pp�WW-#3�n��z�f!�3��JtUW�����[�:��}s!�LHǧ����͆�Etk_��Y��E�L�+�f�L��9wU� �ڻ�}NWʅ�k�S�&K�,+~%����C�X/%5|R�͂E��#Er��ϭN�Eܳ��O[,�DT��:�C!-ҹA(���PJ����b�?�7�G��n�$��Z^��^Y�-�����3�$2s�鶰dCE��^�<�-2{I��VW�B�+.-��NQl�R��(05Ԧ*��N���%��]���r!�H��Q9.��%7C�۝�iDcS�P�/�M��Z`t|��z��$w���U,���d���үm%�U�(��lv�I�o�M�����i�*���mv��<椗�=˸Hv=���2�Es�.,�VC�i�����/����m*��[#�ըu�(�$����2�ƟR�vt�)Xo5�E�J�S����=)S�/�=[��1N4m��k�>�܋���Kb�k>�ơ�z�^d��vZ��j��ɋ�-gk�r!���5y��&�P��+�x�anm4���K�P�AЉ'�]Jt�բ��?CF��Q����6���d0��{�C��0�u^7P��^�9��|f�ێ�[OWk�:+�b<�P�w����-��x�����w
)��ZW�	y�]І��Z� j��Fi��5�a�.RoIHW�_~x:v����H����|L�h!�!L�X��d��i%�1`0k��B"1����r�*��k��� ��y�5�MO;�"�6f���?S�r�L3ė�4� aZ�0�V|`����:�ӊE���BDid�SW}x��F�>�L�~7n_�{L(,����><��.���	e��`QH��c���׬G���.^Ќ�E�+���Iѱ[W`�t=����1�/(�.�ajN�(�R��V���9�h��h�Z��3*#E�]��G`ܟ�j�b�:���@ŧꚟ�����,�G�����~
H�GW�1%�܆��O���҂ѡ�\�G��J�ң�������]������1��p��~�Q�Z(�������7���ʏ�����`�ŭ����X�x�r0�f�!�[��dl��Bn�H�d��~B��)��R��~1Y��4��e�&�ϳ�U�ae�����wF�YָK��m��V��cDʅ����e����~.;����_pp�p�(h������n�Vq�NK�=c6��p>{ևw,�$@���a^,r�����^
����v4�0�ܓ�n_��a^��a���3����㪵v�W���d\�I��D�7�@sg��O�L��v�~����q��L�n,�u�u�K�$$�bd
�k
uQ�it(����tl0$�t�u	\w������ST���6�K{�~��� \p�]���uڔ�0Co��D���G���!��[�0����g����=�����;uh�'^�������M PEx)�[��eF��ccLM`������7ʖ����w����vzFǲ�bsO|y��3'�/1o�չ%�)#nS*S؄��گ��!ƭ[h4�T�h�7'G�p�Asf'���b#���4h��J΢d�.݌}��|�q���){i\�M��@���KL��'\<���G:�Q$P��l��%�{a�s-���n��5Ѓ��<����#��5`6�Wj�(�Py�v��'B�C �������Uƍ�&�kǴ�3���eK���M@_���緤�s��&XW��/m���%��7`do��"���5��;#���&R�$�tg�����~{�!o�-ƹ�48��-9c�܏@Dja~�s��O\�M�J�f̅�Wrn4���,�z�c�����<,�����.ơ����wG=r�6�#�����̸S`����W�����xG�ŔK��2���=(S��=l�v�%�=fj���	uő%���`-l_�5�u��[���p;��??Ò�ȳg>حIzP�_��Ȫl2Ppv#vח9�`�����|ɞ�;N��\d��,Z&W�AM�.�H�aD�i�Ӻbwpi�a$q1[���3���� �M�c��v9�<��ɳ�L�P�G3..�.��w7��Y9�&uІ�g
��C�=@�q��D[7���߁�|ɐ,5x��pٹ��"�/:����-R��EL6�I$Ӭ��7I	�:��8�Rq��<g0U�~�A4��m��b�i+b ����i���EkU�$Wa���R5�*7��xE`��Ay(!����a�'x�?6�����a���	��D�b
�!pb
�Acr�	�*Elb���`�	Rdw�lّ���XJ}(�Ϸ��:v�`�s��c�<������ߟ�utl%�N��Q�Z�w/��-�<v ?�V�9�*�R���>t�{zڅ���(��M��1�~bU� ��o0@O�����a�b}y��fS9�m�/��h�)R�Q'�S#��`�P�	�6��t<f�W���
p�[x���"�s����ն���&�IUWe�'?�=�26^5�my�\G3�I��D�ճ�/@�.��R�x��Y;.3��Zt��\�7��� D1��9|/���-A�G��\-6���7e��"n�����;���kQ�{�u
N!.�G�wA������{���5' �# �����tC���\چ�cm`�.�>����`��)��I�H�!R|��F����9�p,i���R���Y�ǩ���ןtFN>pm8������.�fQl#�'_\�tAu�m�p|0�Xη��$J|�(�Y�/8��&a�Y��Å��P�� o{u~������bKM{4��0v�I���h3&բ�tF|�:���"*�$pPT<�V3�v��*�`h�PP��<�F��fN��lE���jz\י)9A��Æ�ߏY?"ӝR��4�v�	y�N�u��%�FD#�T[C���e>q���m:�(�gI��_
p_ig�u+|(��9m�Ir�=���@���͓����%I�~%O�ѝ�������H."�Y/V5*.(��/rۑ�������e���e�q�Wy��̵�� ��;�lD�n��.	v� �`��9�ӝ��J�́�]�׶�=�Z�tNPS�<Zay'Kr��_��UE��Œ�m��d���8,�T�u�?�[�#��,%D�W�6w��=v��i�s���z�C2TӒ�zYd��P�6-�r=��(��^���9�qA�h( RǂOr.��w<]���Utѷ�1 2~Rw��%0Ʀ�(�%Za���%Pÿ���SiZi��_��F,���f���)̆4��%�	.Y3��j�_� mg��[�|4[�׸>6[�~�5'�S�R�V_��[�'�x����D2^�J�IEvR��[4�$��<����R7ʓX#np�l�')����;]����"Bǡ��0���{,إ����C��d ��C�[R�Hil�֓`��"���E�	y�Z�#�+߲l��5�c�Q��r{���4�.�����y��t����#��f�z�<T��̻]��[�?{]��OW(M�H�=ҍص��Ӝee0�ێb|Ξ�
!��M��Ϛ.�	���/i0��.��{zL���ՒF���+n��J��0#h"hw�ۡB�"gG���O�{P���7��"\c_�sQw������T�c��tk=%�p��|�awG��G�V�Z�=.�ɞ�h��r��pn��R���O��Kۺ�\)apwQ���P�����wH��'����C;�t�{���3ϡ��L��[ 5����KɌȼ���Qd� b������{� �[b������*˘O%wo��9Tq����(ۍq�3�ؤ+��	s�:B�}�3��L1=�2�������>����8��y׶����f�rF�5T.�Ֆ�,�!�zϐ6\&o��yоE��Y%.8Z��)��X��r����%����1�2M�%$Y��4���o��Ik��]��J���[
��<�l4N=�VUrӳ*uˤ%��ԛz����sT���/��p���mT�	����*�X��*�`��Q�q{�F]3�B��,�!N@�XO��Al�:�h1>0چb,�y�@�JXL���GK�ڴ��n���or�c�u۫!by 6�vH��:1��t?�ۉb$��'N��	��ȵXJ�2��f����g��ǂ�}�$������������lx���������/S�-�Mcf�wl����U�u���aR��揾��X�M�dV�ys9�r�x����5H��˵#��C��O���tT�����/���ŏ'��~�	^�f��kRz^=lڏ	�i"�:c2�j�(W�>��N�	[�^h�m��d.�$)v�,�N�ɐW���5������>v���E'�0夰�����/Z�
7\$���`N�$ o8Wsj�	��r���"�b��v�6��n�*Es�p�;_��5�O�;#AK\��^�^�R�N(;�(���V	wa�}be#��s�,����wg�D�{=X�7m�ޘ��WH���eϢ�:�NQ�v���}��~�+�8���W���`�ȋp�+��U~1�0&3C���ߞSEV��Mg苽�ϫHe���i�x�T����g�����1��F�Zӳp��7�L�~�I0��e,Ӱn��cBSb��-1�ii�S���Z�cY���mah��Ë|�&3�ɋ,���q�0��B�)=Z������{��z����C�g�_c�����[�:1eJc�vO��-�����~+;}dpo�d��Fͷpȿ�'�}�aK���^���2��J�|b#摹"�2#lS+�w_�/OFR�O_�-��ؐ�~[Rv3����[�T���uq|��f�\{�}�uj]D8�́�Y�ݻ/��=���CՔl&]�T�g���G8&���f/���p�c~3��ߝP��i�Z��kX�f�Y���*W[�åv�f	����#'H�F^i9��{$L�ͺ���M4!0���t��$�V�j�~��B��^K����z�n��[ʹ`���_/��/�	��3��n�N����^���W����0i�&�o�b�s�[4���K�h���i���oAC�W�>��#���P��	�ry�믍̵���	���/� Y�@�y�Ebڡ�#�}�����C������W���D�bW��aſ���8=@1�8[/�W��Q�ť
@�P��|���EfO&���~�~�㜃*�٠%�{V���
04w�G�K�{Iى��sm/��@`�d	a�Ա%�k:L
Ir]XU=Ξ�.E;��X��T �1�YJ�d@æf�.I�q!;a ��*l��"�ym��6x��3�N�O��?@t!��c��f@�N$���N�RU�+�)�������[�~DW����.az���\�
���Y��r�8��Vlک�O�%���p3��8>����� �9� �F;�:�;/Va�"���(�ud�j�fIN�k�U;t�ILޚ������ZLr��p�UZ==DI�=a��'5�
�W| 6Ϣ��?LP�N�Ur�����
��T��q]�I��]�t:�5./M�Q�z!�g]����-�R��K��>�C��E�6	�e�"��K2���B�HxT��]/�fh�|*b�U5 |�w�C�n�Ft����-[� )<���I�ZC#�`�r����iv���������m�}O�cX���)��Y2C��\�F%��G��c��zxojE(�<�4�-*��r���>�Ĭ�UU�<	xl2�I�f_�P�؄��<Z�}���j��Y�af��Pr�0j6�O�]���a����PpIܹ��Ɏ���մ�X�y<���	l��h���F��+-ݹ�)�*)a�4��ㅂ+Z�rxE��J��&�	�O�yb7ŋ����U)�Y�wZ�&/!����������s��3��AXx�6cʎ�7�� ]�V�VJ\K��j���5�������G�|Y��Ɖ�:u�1�]��%(24h������C=�Nf�̠7.�NL�k�h�h ЖDsJi׿�As�xH|�q�V������]�"�HWww�TU=�}�4=����aǍ7LB�a�ԭu�S� �x�Ӂ攳�;	��h,4�w�m����{{;�P�ä��at�����Ԕ����"U���eÒ/d2�E�-����j�J���W7V�_��]6�iG�}~��L#vO�g陬�t`u�P#����l�)���h�CSC�bD�^L�@��z�Y�쉃����K�I"U��%&h��o)��e-'��;����tԙ^� ��
�M�q��������
��/p�2�_�q�����4~&AKe�t+����W��-z�MX�M)� BI'Y�e!R���M��<u�dz���b�c{��f�LJ�����^�>��],uwx�L�?�̽��#�t.-Ʒ���M�19��e�J��F5::�|�����=�^����0�t��x �S� ��h�y�BmL���C�{��n�^2z>�b]�f8bI�6ՙ��前�c�>��L���!��=�fLS{�)��Ô�L.X;��1���ݐQ%�8[j*���Y�:f~r:@��D�x|YTA����XF���H����n��4, �L��{	Ň�����K��;���6��h�6K�V�q���^O,>�ʗ�E��W#�dt;����V"K$�DŌ��[��%6�Z������D�DLn
�Ju�����6�;~
��w��~�[�b�Tj���ˀH������E ���B䱎�И��E�п:	�z�Z�>"I��;"*�m�t��2�m'~ ���
�1�pk������B:��͔���J!���sH�v��b��/�U>�! �d�!o:r]���yh�-}�r�\�w�(}���	�Հ�>��X�fF��M8A��2�q\�M�l?䲸7�3���h����~Q�tO۰J�GHiY�]���A74�W�����O�2�QG�63_q�j���x����#�g%��?�uKw�k��P��9CBd2�ZF����\��~Ep�|T_����(����n��Z�������-���-bZc�{�I����4b �s�+�z���q�`d�*S�	mM+�h��U��Edh5�C|��B+��!ߣ�,j|�@@ǥ`y���Պ��b}�����[��+X��o�43�9q���Ld�-�D%/[���%AE��,ve��a .����&b�q��v��������g�^%��Oh��Ě,��������RO�m^
#d�<�V+oX�57�D���ea������i�k�����:���ӗ��z�^�O�H�0V7�K3]����4?Z;a�O�	�O���n���]�l��bFAc���c�%�!��G���_��گ�=B���AZ����X`��]�-��5��5Nc��O�����} -C�F;��ټ"�y���py_�}I��G�-�,���k&f��K^�2cm����eF��0�j����'{R�3�����Ȼ>����8��d��J�G��Ȱ��.g����%`D�<�O1��u-@O�C2�����@�ύ��0Z����Nqx�MLMF�[XY�4@`�1�,n���݂oq�<�>U���K�$��S�gU���5��l�?�+-MH��|��I��ϔB t�B���7�4خ�3W�)ogB�S0=V珠׼/H���	C(���G��Ft��4�|�S��NIn�u)Ihck�D���١eC�s��>����������;��RhIK��K;�F�zY�=��?	�m��3];��K���}ˋ_z�#�� ݋�\�C�d�z�o��Xj���UX}_C5I�.�8��}��1�h�Sݥ�:�!~�h�a*d"><)�'�k�r)}�5UV1Xu��1��az�r�VX���`�9*�P0���Z�̉���dUr�X��猳�Y;8l������(=��"�m��i9ɘ����&�&V[���D��=$���	�X�"�OJ��O���ڞvQIvZW���C<�g�^�e�?w>9.I�op>����������X�PbTKZ"������m�!bD��=���𧮿g#�N�~D��O���(ۗ@���8�T����&_����4��?ZԻ��V�Gҝr�9+�zz���"�@�Ik9z�R�v��09�6Y�d��(0�{��|2�Aa%���f��� ����@��*9R��2,W���3�k�,�ȱn(��i�u�?�8D~�;��h�5�M������ 2��9x��#Y_�ݫ��[Zh�?�9?��5�!N(1��{ޫՊ�s����}��Oܺy��g ��S�T:�|�ʣ�B9�~׀�!Y��*�ӳ�i�j�����m�E�sh
6����ow�U;��88�-��GY[��������ƈA��fq�`M]�4�Åd"C3�w�ֆ�v�I5����ur0� ,�j��_�;0].�I�a��J��,�E�������_%�|8P@��#ʉ)[���J�u-�4�0Yn��z�����jlۃ�CM��c��+��-�%_tjl�[ �KV����e�{䨁�����	" �F1��֐#!i�?uF����E����%_�:��_Ն�_���|t6QP���-`fY�G��v���ů�`tSӔ�f�q�1���3���0/ī���R�l�|��xA����B���b����jWß����C���L
�@w���P�B����@3X�k�X�]�x�$�ͬ'H�i�����5AZ��H�lC�ET|Pk_�z�Ӵ.F�ӼKT�3+8��h��Tv��W���h���>�P6��:@!A���w��N��JL��^�*��P�AbJ���'t:M�r�Ă���b�����6"�{j]Ac)\:����Ģ'T,T�����
<,��!=�"�(�0�dO���������%��D�ѧ�vzYj�?�`n��F[O�ܭ~���o&�������Q6���.͕��P�ߋ��J�t���˻(�>�5oz��"(�~��?�����ך���@*��7^څm\D�c:��C� Qe\���ēR��È0�֣����B��k+]��M�L����C�.��M�I?��ЗMϗ=�+�ɪ�Q�>�0
`�}�U�% �n�!Q�vEn����Ti5��,��A����~r�ř���G�+5�pO���t�M䶊����^��r�GX��,���-b�n��'�B�O��%L6y[ƫ"��zb����n�Ww�N�ߊ��n���Bs����Z��d|�������k�B_!�Ұ!��ˮ~�]>�]���F�-�!k��?�Jѕ8�|̡�<5Q*c��B=Os�K��ӝ�E  �*7�1k��`V��K�uf�֔��6�8���������S܏8v���K��9��Fl��Z�\��7��1�,?�?�E��"Ťߖ~��FY�;o�l<)4�/
���ط�*JF��i���#r��=P,�����4jg���qm�>��C��W���~G
�?�>-};���w5�s�U���4'1�:
Cp�tei;&�y��M_�;Eh�|UZ���pPV��j:-̈�퉃*�����Z�KRW��!�=������-��F�H�U�%�r�<�����Lxy��s'F�**�dR)N�����Z�[�	?