��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�YM�C����ion�W#a=9�-��R����R"��@��7x����\z+�6�ۍL���>c6-�7ݡ�;�F�Þ2�[	_�R{����p��,o�"2,-G_cD��ç=L��C��������>����1-�4:���M��;�`b͈ϧ�4j�wh٘����b�DTʶqR�)dݗ��ѱ����`8�\��أ��/�7��c��\��0j�.xD6'јN���n7��gqfl�w{��]⒠��:̅M����K��$���X�QE]�cAï���`�ׅ������}�1�{�����D�AS0��Ml�����>=�|A<���C����I2�>��b�=�e�7Tc���Ό�#�ю=P�^u�_,l3��.�PO˪a�w�ȹg�O��;��F�V\7;��:pv��:�8��E�����֫ƪvy,���tl0�3��M�'P������A�+ �Q3�P҈����ND�[q���(>VC�u�/�˥d�T�h
�&��fs�#��ǂ�uz�[�~�8TF��!�BQߴ��&�&���N�^/�Hl~�������n&G"f�<�h2��2Ǽ��|�b����N�3�i-�6,�m��U������������vqHo�7h�����.Q�,��=�J���}Rw��QѼ-� ^��p_&��o��O�06�EB�ƿ�3�!��cSh�м����j�M���S�SJkk,`�"_ZK�Gѕ_�ۅV��"1�@�e�|�Z��F�����<F���'jȄ������0)m̰V�_����oi�R���i�
�l��u�����̝�~!�	����� ݦk1}�E\Pf���%����G�4�@h�~;��t#Rgp4�.���$�U��T����<�h09��1�g�BV�X�Dۢ��Fc!���r�e)_�$Q�=u Q4n���`J���GZVƓNM�>j'0�'��@��~ yh������ޏ�RD�oV�oQ`BH�K�
��a�� (9��b\+��B������rx/�b�5kъ}�2�P�!�<Op��#,�O^Gz�n��0Q��I	�V��֕������+������)��W�Z�~ԤG��[���f�[N6��ZӁ׆:0���ڃ���TQ�.
����8 ����O��d���f�b�%k�\��l^��t�n2��i\�Y�(,0��I58:���,��{�e��%)_���(��x�w��Sq���[qNm�kX&��?�Q%�~R�}�'�&C�+-�E=����v�h=4�d�VĐ��Tv,��J�Vu�ǐ���U[�u�O�	h�Ǚ�i�N��%AUC�5!��i���z��kx�x�U1�/��T�R"a������W�2�	+%�>��`6)�9/�mXǏ4j�Md��+X6��T���\�ٓso3j+�0� ���rӣNCڸ�V
r8c���.k�m2�QI'���/��8>�''ӾT�&��~95�X�T>�*P�2��6��Iş�P3|����ʖ?��F��i"i�E,ƶGJ3񣻆H� s�OR/���KL�P�8�2��7C�z��E����ݽ!?��?��*�-w�&,O���t�X�.�E�z�4\F ��52�->�DC~�P{��;���x JG�B�8�I�����ϱ>�vn/��Y,�W.�;�`z�	��������K²u7��د���n��Meͯc���[�Yv����>>��:s�T<�|��;�ec�&����W砳��/�~�Q�I�ݵ�Ε���6�#I���R%de��?eEc�p����9�o���ͫm�A̳t�x��0>��M�DBi�*Y>I�8y�������J�����F�K!%Yx��e�ɰݢ$�DԺDmϲO��X�ۃ`�s�2�} ���,8��e8��s�����[w��\U�S{��O���s�}�;W9F���U��w��;H�� Ą��]�}�z\A�Í�^c5(�9q�a�����c�Lt���ϙ���>.��0(x�(dC��>���P�C�(���8�q���pm�QոodK�����񴤙��ܲ_�F#�