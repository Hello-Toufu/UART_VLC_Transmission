��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��v�N�쪈��%���ieLF���z����$O�� �I?�r胬���TeUͷ���ϴ�I�'O(�y��jEr����د��6�P��y���1K�\�4ۜ�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�i�8����!ׇ��,		���\*�"QF����iB>��r,������ADҩ���'���a(D��`0�����Z2��F�X�ů�ѽe�&�-�I�C�ER�t&s~���\(�@�����

�f��0�Ok|�f���X�3��GS�H\ܫ ���N��5�Gސ�#�V��0޽$�_-Q\��c��_&��Z�ׯ����H*%���s4y�_��n�c������۟�-D�l��U���닚a�؝c$NI��%�c�Q�N�ՠ�<=)4��K@���g���ߗ�Y��u�{�����,��*�Sܤ����;��\��W	����5�]���9|<�Ҍ�]@�`\��]�ز-v;���&����>2K�ޞ�hb^G��r��/Ru@,�T�����we�8���&�y�K�H]V�X0����l#���}$Ѻv��)�f����R=��	ѳ�1BW�m�|Z�<~ڣs��_i�w�
B|��+xW� ̓FF�\kZl֏�F)7)F1~>�Y$.�{���{���z/QzAi/�Q��P~oҗu�s�D�}ߐݶ���=��?�I⦟���'�����6r,;!�-? t�R�?���rQ%Qc�3y�m=�?�Vnߦnd݆;t����h�1�B	��u� .�2W���b����Tv��`{+~#�݀R��3m������4�YM���z*�Lp`�C,�xDgR�6�حi�C�x��Ԯ��뱬�e�F�� �Lcv�ii�JaݹS�����y����̧ye�q�:���� �g�i�/�����Ñ�z�U�\l�ۯ}�[��k���f��*��M��K�a했si҃iG�m�^"����7�A���X���m�!��*��ʷ��G��������f����:t�����uC:����KlߤPO�8�>W��i�ɜ�'�F|�C�����iC}j���5K�������0����/�8�m�o���O����H��%�C~Y���#���8��!D��VI5����A9�.d���)h��|86�]�;;���*8�s�ܬ%KR�B�WDw�[�茛=�:���F�GF�y��K�rp�۲�"L�]t��p��wħ\iD����=�P�k/.h����x���Kiu��@����Z`~\Q���R��٩ݯ:cf
O���L3A���<�_
��;4��꞉_�U� �,������p8��F֍~G��]���b9�w���9�L�Zn�
)o��Jh.C����T���1� O{ywH��R���( ��R�C�#øDr"��n���Ew�Z1�9Z�"��n	����>X<P]��!l���N�@���Ȳ����ZB��t��Ck��4I����Pl˔��4��Yj�8%��=��W|l	���!h:�#�1�?��<#�#T7pO�����Q��5