��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��P��=:� ����(�)3�� 5����l]0�ك[�Y�qޡ�(���fZ��#b�}a�3�
>cO��o�LW��4�C���(C��&{��"�v11#/I�&�)�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_Kq�n��Xs��P1�7�.G��H&k�U�mJ�	�(�1�	'C�2�\�gJ� �a,z,��mi�����.��n;�"o����->�YH�^���_Z���p�oY'e��¯�`Fz�`ʻ�*�R)H�qq!��M����â��x�m��yh4�U�x���V�D�\m8��Lğ�]��(�AVF�+���q��c���|�2(�>�b!(9�14�8;���]
�vL�;�T9ƃ�܂��^A��A��tY�� �mn�t�m�D�د��Vk�� +�e4K�j���B��I6���3�[P$7�1�\_�R.�j���6�����c����>�"u�p�����Z%�L�7�?U�9n��W_��*W"��;<0%�ɢ�$�g�)n�����u��������R-ç!��e}$N-�%5��%F�\��}=���b��
�k(%�b|+���LXc�2�v�?�������b�s�o��Ii��+�"5t����|�q~����lj��E���8>-V�t�ط�gM?�S��w�bʀ���Kf�Z��:|s�/w'}�}��@H��hr��c!�������XB�Ƌ�
N�3O������� |��|Ӄ�m/ .�2�h��h���5!��ɘ�s�éFW&�ݟ��T����馫��p]20(�(G�W���Ը	��	0�G
��(�hH	�b����f=�s
:n�Hix{!�T��i��^F��,|��"�vF��Ã%A\�	5��&m�����8�ʻ <΢���/Y�5L��Kن=���⚉L�[)�lʬ<K�d��F�̼0g Y��H��U�MBh1��_{�O˦T����Q�M�@<1�2���
�O���?R�R���hk3/a��P�ˤ���+�/	Tn��bs����HW�7!�~K��C�2^�5�´�}�Jo0'NSl�����������w�/��Y�=����;,a�F�0O��l`SR�%�T��;.A,�9��Y�{Lj� '�D��ak @��!��>����"Sz��0�34�6�� ��1�~ڒ��bY�i��7(�W ��F؍��()-�E�8�`0�IbT9����JO[Q��0�L��~�>�%����t>�{���V�EJ�H%'T^z�j������Q�fv�g�'jYge�E$��w[�M��
�A�F�&��hI�\͗tT<�Et��Y��g��7؈2L�Z(n�k�T,�.P�lo�5�E#VIk��Mx:@_t��H05�mz�iAAY���dj�<�\:�17ez�������8qud�
q�}��V	�l�f{~��Y��z���h���@�fM�q�D�����w�)"�1����K�[��W��`���`6����k�}J��<P�yO F��Q&%��[�t��9�2�"�Xx�q�И8&�&Qk��FW��O���'з�+%�/�e2����/gP�J��.��.�N�|]\#�����$o���<~�'؝w1ohO\�1*m�6ǩ:�o��&S�.ՙ ���X��}��?�1�ל$Yi��Y_�{�iU{�����­��d���O��{��)i�;�t����Tw2�tB��5�o�w)���Ʋ#�	��\�x��E��.����l�f�(��y�ˀeO����	�%�_q�J�>D���wO7����<��fm�r*�����)Du���10[u��&�bė��/e��		t	_�Z��յ)�����ǂa��-�'*jM�3
��a��}�������k��2z{�J�0�Ӄ183�NP��p�ʡx�	�g/X��t�lN�+�%(+KhO��j�buտ���8�7�#�0k�xi����ӋG�5��	#}v'��'G�R��VP*�H̴J�h'�?R��ᮾ��RU�6}�%?��Р2�Gv��f�vFy7K�S�/_GhO�\a�ܰT�rH���(��� G�D븊����f�B^���o�</��y��9BV\�!�w��γ���t<"�~>,:����aПx�$�tJ���G�T�?ND+�Օwf�ǭM�t�O^fw�@&:���~�V`;���h}^��?�ғc��SJ�_'�rV�z��}�![���#m��+��i>ծ-�߮u�o�b&��K���-V���q��~�#����2��0T&���l�6
6�;A!h��ɟl��A��^PY�+��е���]�<�E��v�ެZ1<2I4V0ٲ��t�[>��k���~�f�E?�#�=��9�g�#���|�)���|�<�"	���+��H��d�Ӄ6��>g h��o���@_�'^3���t���JI� �M��p�,�r�7��1$�m�B,6� e�td��7#�Y�r6b�O]�N���*$(��X����_��^���y�>�AkV��Ԏ��C�u�ڙ
C'�2��~Qq�o��`�$w�G���0��R��٢et�]�2QS�'K
�\X�[!Ygl��Y��l۲N������J({�bL	U��aM�Y�`�q�bM鶓7�K ��Fa�.(uaW`t�ޠ���et�_�D�xt��֧�Feݷ����ْ�墢F�}ָ��cB�����l+�x��G:׾K��n�M�0n����� �)�X�H��W%Jc�����y1�W���k�V�h
.���	wFYJhD���Mv�3�ʜ�
=O�t�L��R��E�hQ�^�s߼6�N�tt���G�6�5�8f`T���Ԑ�{M����f�#��SeO�J{��[�
�nd[���LiH���.�n�L����t��څ��L#��U�KV&T�B���0Jzu����