��/  B!�;}FG��[]x� ��F"��ͽ<�鵧�$�u(��6�X �=>�$��K���<��~�Wdap��L|���8���,���M 8q�T=�j��<�0!�J,���6xR�g���b�o��M��,��C��tg���M�90y٨8�9u��ț7�K���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�?u G���r�bbd�a)��g3ý�]�mv�e2¿�f�N�dv��G~�nu�[vsd�w��<��붦HYH���ܢ��dO"��S��������t˜˺�����?I�t&���V�+���i��A06$�*�!��	��?�=u달^���  �eKDm <���������Whs��*(T�n8��C�q<��}\�_L��]��҅x�� ��	�*����E����,��ǜ�.�j��$��e����8�z!��D��ϣ٠:���ɚ9`�7�j�a,�!�]p&���]���U��(e~ꁃ4��Z٫��u(DL��>'�r����Qg���8�� ��{[I�.Z�|�Γ��R��lZr���ƛ��aSKYR�Eu��f{�P�~���}*�F��w�?����u�gI����UNK�H0�nw�������	G�OR$�9F4��,?fNM)�](���+yf��oN���d��m ���,I��R0�g-�vK�Br�S/u�f��q�x��?�v�j�����|�Mج��U��g����#�n����CG��-�p'X��Q��rH�R~���$���8�v0u^1�nr%��n;_ߊH]<q��1��aṞ�"��l7�-,=��V�]�,�#�rԿ�,��?���< Y��%Rq�փ'$c��g�1�Y��	��N{���S҅Z�֖DT���ܒ�����Ip٦��bzAB���S�U���p������TjEf�����Ċ�ha\��T�ȗ2}7F�ɱ�X��x�=A;�ַ~ubr���/�D�7<�ŧ�f��_7���1A��x厭[�I�F�N�R�*����NB��/?�ԚGǡ��^ ��%�)�w �;��w�)���a�ͼ���w��U;�i
�T]�eM���&��~�I��#{�מF��N�c40�H+��́(&w��,8k�=�z���i3B����|�?��N���M��@�/H�=�\-	�q��0���S���[*��eTj�dBMV�p.{ݫ�n�>'���;ޘ����M�1�������4"`7�[?6?*��:�*�(lZ�������ﲿ��c�Y�N]��f�w�������f>������0��sNثP\GP[��ҵ[���%P��Bp��/��Zo3��x��̸V�(>+�B���Z�/%ma��z��FK,�_�	�z_���`8C�� �t�f �N�.}���;�K?�"袉�8�4�>�1R�RI�r$r�ڌb2&�葼�\��F��-l�q� ��Z�Wqß�'SS`�2�:_��������)=,|�NlJ�/�'J���������P�U���z�*׳;?���3��s��Mɤ��?��IW�~Fr�(ȣ�%B՘R���Q��}�gO+:�=x]���nV�_��ϲs�����'Qs�!d� WO�	�7z&)�`�@ș��畮e��b���h���h(mb;lS}.��e
ѣ��-MK�Q�u�wt�'	��n/���aP/�a���*��4a����������=K�Z�O�6�!J*^f�=���W�2�+v�Ib�P(·�E����R�>0���"�c��PȂ��_�l�˷	Ճ�ǘY\o{{jP|�&�����9� R�do�;y )�!-.C-�)����K��dÛ���r�~H]ߏ�	ΚA��t��	�}/kfGX�J���wcУ�cZ��d4p�);A3h�xDF�`̰����e��-ݺ:��H��:Wg؛e�Rbn�ݻ|4���axV�EY�3{��OM��/W�T���!y�a��џ���ۍ�>H te�n.)~`V�Ȩ���W���Bہ$��qf[j���ߗ�>q�{vE�������0(Q�GJmŧr��8�Gyf�����K���1�ŋ�!�`�����*�N�@���2�����n�\�j�ԧ�}1�X�� ��w@�o
q�T�U�u�P�ӓ/R���Tf���]�v?| R�gq���<G��]�@kyn�Lo���rR`{�gD��� �"�]��"����D�/?�HaC�\���Z@����4�_P��ۅ%�;�[?C��h۷LG�*,��]�N���-�!^���Z��*ơ?g5(I/ ������f�b�G{D��ᙉ ����RK⻆7���W��4��ݨ?�!U$R��I�$VvH��F�T��AF�Ny< �,�U����A=
��]v!B�;�3����N�j�1����G�񃂷.��z�EqA�o�\��R͕Iщ���&qQxqݿ����\e���{�|] 2������Y���G�El���iO�����s��;��<f;Me&�k����{o�L�+-��D0�N|�Z������b��*���i��|ĩ��*;� "].<�?@�RhWѸ<;b����f*~[x�s����qނWm*Y\����ZΒ��7��[�����q����Q�
�V!ﰦ��sh�F��Ơ�%��>`�l�SQ-��H|L)c;�U �����r����Dt��h�@��d#�xT&3�|�����q*͚�r����Ǥ6��l���6��^9-�=���1��<b=30bN��2�����c��*U1Ͱ�6����*60�T��UvF��������A=t��бMK�=	�?��] ���7uU[�S��zR��0X�ܺ��R��וlwP����S��It�I�,�fP�
�e֮>�"�C����Jn�W�q��۱tӥ�����"շ�-�9��k��iJ�U-N�s�fp��߃��N
�qDZ����܃�3� �ˤ��P,�%}3��v�sN�	��.r��n��l��8�W�O�\��eٴ�Mc`�9�J&X�~�,�;o�����7kd��0�<�R!b�/���`�Z$�v��?Ր_{��ޛHc����������# ��Z���0c�:�撶��R������En�phJ�����kjQ��CQ�s����X�ӟ� " �5��9�O��ל7Zp�>�����d�c+R�
8�s"+�d�Hzw}1�D�����!�����'�@J��k�o��
|=c��	���(\x	�y �k^�,~��|���/7��K�q}���q��Zr�}IL��7.�[��.��n#��`��YklX��8�\<E4ڀ�,˴���㭞�h�(i|�&�����
2f�Y���^b�i�YL!��W�ѧ=q�fz�~_�4B�.�Q*��q?H2��0H��~�"��}Փ����͙���Nkl("�A7���@�<9�&`q~���\w{��I�;���������񩽲:�kz{����k%��\��ɕ-ex*|.�=� �
���ق4��Fk�����H]��_|��I��W�dj�L�̟�G�0A�N�8'��f�&aq����	l�_��l�s�t�n?�y�F	"�st�� ����*��.�.�s9�bH����R�e�g[`��R�������W������AhO���- 40/���N�a�8W�!��~-v�B�-��<U^�Cco�߂nf��L���#�]���7�N�Ye���6��ڜNf�G�Z,ߏ ����Y��̚K>di�{ѱ��#�����<H'88|��񕜚���u#��x�u�ef��o@�k��K���+��9�b�̊'�C�� r%���^����q�cQ��U3����gXr4%��)�"lHf�_��_?�0���d�a�-���T��?�#�V�W�n\�kk�F��<�f�TXƝ\^(? {�-m�a1�����7�[c��[��Bo��u}P;Z�>���/[Y�[!vS)dh��OM���耽�-~p��jMȬ�"3� C�PYx�s���V*���B!�v�TY�ơP�Ts��q�y�~9ҁg�g~tG�ߞ���DF��Ĝ�F%S�|�]����>7��S�q���1`��Ub�n��r�� dk>s��:����c%���U����wCZ��"s^�$<+�N�rIl#�)�V�b���jE�m�$|�ɑa���}T�7PҢ#tx}��!���N^�R;��Y����2�{]�"���P����_�1j�Έ[�;և�_��s�V�ۃ:��C��l�۝Jbq��u_��~^۾�ɓs�����ƪeB�۔�����)�R�M�D�&\2��Х��*DA=�&�ha"�K�Tg�P��a&����;��weASF�,��2����k`h��	*WA.|�xQ؋U�p����֞
LW������+*`b�gq�u�������.Hu�`-�s(��8͝�`�ѡ�������Hb�P�q�ãW��W����4~�K��&�� �9�O0Pp�]�z���@Qd�0��Kdy9ay�^��;Ld�Hh���R=�g)���^�� ��=!7gg�? 7��S#�EFR�u-���k ~��1�O��Qj��v�V�	�,C���:���GE�:�<�8� vs�>���f�L*�#-=�{�|<���޻pe�	�-D�h)���߇�,��n)��'?IY��scu3:L��轆N��b��J$�N5��?��4�� G�L1�}m]�.Nt����l�'�o��3U���I�G�Ҩ�K���Ɣ��2R�.��E3�ce����9K�%%�@+��ej�u��Ȯ��[I瓍!��L�n`w��\�����b%'a�ɛ��U!)=�mS��s��Ơg���W6�z�^���d�������6��]�|�U�1�h���a��j��H=k��%����=�Jm-�cy oi������g}Xt��A�*ꡚ��ՊQ+ .��"O�f�s���?5O�K?C^uUa�`����x�Ћ!�����\�Uv��;�wW�ʵ$s�+�6�&Ir)~t;w�����T��� �߳a���Nv�|�4���'8jW�ۣ��̟	I���V�R�߀,%�{�2��ȡ�@�X�<���ynp��!���s824��I+2�=�.E@��"��. �.��0�Ҟܸ� r��������P��ԁ��)4���0��ia �����n]T�j �A��?ߤOʇU˙ɓ�/i�Pj�W4�����C4�R��c��S�\�)��δ�N4�-9
�/~Tּ���k�� q��$ȪFy�5���o�rѤ�Y&cDx����Vd�����$C�hdC�7�ۜy/���X�z��^��x�g�B��3�&��^�ǞT�� ��O��ʊ��U�����]�X+ݡ@EJ���񿘁o�ꁠ��>�V
gÆ��h��@$����V�ŝP�Z4�;������7����|c()�@����"㌻Pbټ��۶��jԮܩr�9�x��O"���J�je���%��@��I�nU�R���D�[�e	��
d�e�-����n�`����L��_9��
��F�� .�a� ��lOI�ߴM+ޢK�%-��v
����������>%4�v�������I�X�5�~]bF���KHǓg<�w��g��=bY9�]���&@��:��x��"R���w�(&c5T'Gy����=-4��WЏ������/�)N���� !]��u6Ϲul���B�w��%�Nx'�_/���} FN���)G?l�)��)��P�+ׄ����n'�<�^hw�h�iX�_�A��)A``�FSkY��h�A��@w4�\�Q�W����
�;��"Da1�Vq`{g��y�s�/�P��n*sX��!k����1ˌ�4�`��$������ARi��+��S�I]��|B�,�7vr�*3x���9� y糧~�O\�_{H���!,�Y��9`�a���l���Nf?2�J[T����8)�u7�(�%��ߑ��7�?�4�J��4�����7E׋�бz�x�.�|=�X���	ҸQxHr��t\���r�%�<�R�l�9	����,Ph�p���eUr4�Jz�9�2eu��g�Ӯ~U���㰟g����&���>���tBRY�²��/�����/Y������e�����ه�TL�D���H���zR��#`�Kw�a��M:f��ew��D����,�Z8r�q��f��j� �6�q�L�����F9�nޙ,���3�[���k�+g�T��u��	��[|���Y�au�F��_��m��� ��P���8C�N�� է�0���6v�
@��S���B��1�cd0M�X.�򧝟�ߊ^+���vf~�nx��L�nlT��ub�.�@8I��ڠ� �VA.F�N�wě$_�Ԡ�x�����ITky������ 
�9h��4�:O1p�g9�G���Y<��I�@]�]K�YӬ�h�AE���^�i���t<��Q�rŐ��򠆜x�k�W����u?=�}�������/�S��3d��	���6.O���!�>��K��UqA�+���,���1�Ilt����gPG�έY���	�qZ��(	϶�1�B�F-^��F%�XOV�U���x�R ��P���oL�i�`���w��`6�٨������Ԅ<��В�{�R�
�X�'_�h���3�}0}&����a�Fu
�t��:ۡ�"��� ��z����$�~Y��󳃮�qL�a�E�= ���k��3��3��Ŷt���P#\/f��λ�n���:����r\���<���Ⱞ��*}�`B�}M+�Kqx;�l�;Nze:q�m#N�)`ġ-��^"|�0�L9֚2��p�����i�C%zk���+���-���+D����3�X9W��^��H�H�����ҿ���U�EëO�TMx�-:2!��,�����i������

�AR(���͠Klլ��!d�$�P�
¡]2��r�+��s�����Q�蜘ԏg�&�:L<�6
'�Z��z�A޻�к�m��D�����eo3{��f��Jq�bChᛴvM&�G�pl�dy����m���$vU�k$Y�^���W�U0�CP�}�/^�DKK��Y�Y2YЖ���`����2�C�a*=T�ئQ�2W�c��~'��6�*�̑�B��B��ծ�;��؊�8I	Bp�����IA��y��G�w	o�C
��ڒo���@ ��i[�d�_���C~ӗ�y�L���-����K��9K���O��ߡQ��s[6�\�M�H�S�L��PÚ�yoeq�;n�o6)��b��B:����My��.g����C�1"?����TN�D��\�H�*���ɚU5�M�2"*��DQ'q`�ov~12P��^*fрf�dO��(��C�Ge�]�L?B��4�{D�#P2[g���3\LG�L�S�Z��:`>�� ��\�?�c�wja=&�KO�eB]W*���v���n�'��'�'�9+�-�Kh�͓5G�KQn7�9^�1Bh.�zҍk�C��ڿ섾���^�GN�y6ֈH�O��~nJ�O1\k=�h�Q�DB��~գX�m|f9�\j=��Vlf�*���N@��f[�I���ky>�۾O	2�(�,wEF�F�����`4 H-ʝ
pm��ʻS��"�Cɿ~M{k����]�:b��?n|����3f�Ӆ�a���p�s�K8mi���6�=�mr��&�m���q��WW������Uf��r�i�MBX�X?���}�V�Y�l}/|vyfw��-t*?z^/+���E��[��r˖rq�@��>���X�?���������g�ͺ [�Z��AP�y���kM��X�wɾ�^\7��
n-ԧ. �Z��Q�oz� �k&�+�jd���W,�!�c��mbN�\ܵ.��Y�'8���%�z��p&�6��R�,z��ms�J�S�d> �����f��y��:�}Z���-wy4�q�5Z�#�S*U+�U�y�;�m;�'�VD�I2�Pb����  Z[ˌeL���p�����ύ���c@��g�T�q���H`������p�VL_�G4� ��D�Nq1�n)�G�H��^p����-{�@M|-uI����YYZ�(�?�:���h�"��16�\Y�go"���0,�R�)͹f�T��0��p�?�̩,3���4�s{7%ˠ�7i����TɈZ�wB���Ҙb u�p���4�>S�w���Ѐ���'x��=�3Co+Z���қ��YE����
��˖'�F�|O��zն/u<Hn����?�THa���h��VS����F��C�δ*���M��&o����@6����v3�D�M&=�1�{:h��*0��q&6�����k��G��/�],��͈iΕ~'P�I)|5o�1�_��ˀg�ֻ�>�U{\nУ��uQ�_,�����2��[ +|	{5�0�|�//��p��V�������a�r*/�y�5���sD�x�o_���5t���ձ�	��K6��_#��Gz�e�S�<my��*���K��˕+}1K2<
-��#��dZ�*��nA�]�)�r�A_�Ҏ�>��}1�Z���~R}Omm2�
�t�y�-R�t)�ũ��@�c�ś�6T%��y�8���v�,}�-_!�1�D��&:�w/7�<dci�HiL�pKeK�ӢI���~�������󻜋>j����l�9ͨ�PL��3,��Xv��Ȱ
��J�ѼzK���u�E����UC(_�W� ,�9��;#�O@��q8׃W;w�o0)j��m&�u�h���;�����|}	O����A��z��,�\G�,��dÝѺ���)�z�+���#��r�xLa��ns�ш��	�1j�^��_r������DG��00�W�|F}r]4�E��v͹���,Į�CV�O�����y�! �Q�o@K8,�\\0QpB��QD8����/�SRzx�?�J�0z`���4�5�G�T$���#�Q��;H��:$\�!��]Nџ����Y䑅0��z�]M�.9|���bŜ,W�<1��(��Mj���j��l��%,;y�ԫ5�Pb�}alg�,t��P_�>�)�p��'C�+3�*l@ ~N�#�g�<a@���_�Zs�;�ro�rW�s���^ҽ����؞լ��IH*֐�@�FN0�����+�Wv�������0�����O����.P�@e����l
�q�RE�AT�C�?�C�L����g�y�6�q!v�UQ�c �OQ`x�3o�ǐ��֝f�d�$�-6b �'�V�D����F��eT�m��5�|,#���a��� �w�9Oژh\�?msI2����i�Ydo����8<�M���l�<�hS4;�J�78uo��l.8��Tqh�{�l�s����WX�8�9��9t�6�d��1�r�_�wG���׻�TDb-�Em? ���ތ����4yy����+���c�#���M=�5�����x^���Ӌ�c��7S@Y�y��W�q�v�sȇ��
��!NMq���\ ��y�������� �p	���M3qD�҇�3�O+&�������z�_1p53��F�[����uϿ���0]	~� ��~��B"�ǩ�����,BWב�!���a�4m]�!	#J�e�B�Y���t�v��x�a�L����}�"�ٟ�)#n�m�P�+�*q���5(ja����;�	Ğ�q����{���^Q@Tw>���z��:�\��7�/�3�}��(3/�~T���Z�r@�κ%�q�^���:�G�23}��1�c��S����i��&,��A�;���ܣ;M�Fv�wt:HUe�P��3[g0�AY:6�/�hP�H��M:u�sp�>RH�<���M��9�kc]:{ Xچd��0"�C��l�\�3`�.�nq��l�jT����s�ڿ�j�������	VZ#Ã3��k����c��@Y�%��%�R���?�Y����|��d���[�,��'&�5&2eO��<Ż������ꈈ�D�'���/Αn�n��'>ݠ�#I���<E�����M�Q��F0K��e�c���*��8��@��,�,���L>`�KUE�Q�a;�a���x*V�%�/�i�!��E�ӂ-K�8jH�J�ZP�����j'���~�Y�p��'$&��-r^Yu�؈�L�!�R��y�$�*$�#ذ��:�`Z�7�n��&]`�~H�Fxv;��l7��g>���~�nү�{N�2�l��wُ��yv�؄��"Wjj�7�iB�7�V���Y��<�e-���BJk0��@F���tA�3'2Ȩ=[�.he�R��!�K��4N
Yh�H^���td���x���?��h�ϥ\�E�\,
8�C��#l�-q�	���Ǯ~�N�ZW����IN6��	����퉯���B�t�IS��'Buf��X��ւ�!�Ҡh�p�����A^���Lϣ�l*�G���C��\N'*;e��m�{���
+R�o_5R�ܙ,�g鍲�J�w1���L��6d�ĺsy���?*���풃\ݷ݇-�n��Kxcyj��/��W~h�4u����K�%[��^�˧�R�c�~�Dˢ+�d�D�ZEf�A'��9E�5<�����[�c��}&=�a8W�����(]�c�8P�ߓ�������r��CQU��1�H90w�F�3�gŁ�O������O�(�������^QJ�C������z�jvA�b��RkB�[ʹ^-t�)�\�u ����z{��є}�w��sK I����x���[\Q�c����I����)=̒�ay�ܺ�F��R�$PA����ؙ}ˠR@�N]�t�+@4w0�7_)�T��"n�A�� ��nz��I��EJ'�i�
�[S���&�`7J����.��g��PI���%�ud�q�ЊBᖸ�����I"�s8���N�݇�E3W��~:�V��ҵ�^IYLe�By7��H�K�2�~�ש���Ћ���x��r�̑�l���=Ӧ�p�P��Վ��/j�n��#�0��ײ��-���8�|�w�!���Af4;��a�m�""����hT�Yw�bU�v�〨�_��}�U�V�t��j:&�`[Xj�>�~���вU�W��<A/R,��vd���L�aJ(w��ȷ�p�e	d�=�X�<��W���F���Iã��2c#X1Z��҈����ֳ`�X��;�_���� ��vS���]e-?�UO��礈%�	�o
H�>[h���u�8�Bu>�sK��	�����^�n����&昺��jV����bb���!�qS���\�G�r��c���S���%�������Tdװ�i~�|�3��Ԥz`�us�mq�!�4F�tjZ�df}�-�]�N���7�,Uķ 1��Y����y ���D� ;�%��a2h/�0��K�>IBciin-�u�w*�`���	�qM$ <�%�����BJ��ڕ�v�4��d<�*���� y�4�G gy�	�A��h4�#��ܤ���?�Pxh���5��Y �9S����d ���L	u��ra���R���z�'�%���&�#\��'4�%����2� H&�kz\�k�X��_؋ҧ��o�z[z,�E�ع@И��^�y�$�ަ7hۆ�����O�~��ur�����c�^�|��ϭ�ݶ��G"Ӿ�w���Pu�m���՘�%'��V�i�f2az��",��3��y��XY4�T�\�z����˭���el>ㅈ�j�1�Z��#��D�K�ڊjz�(��f�$h�/�ʼ�ጌ�f�c
�����U�>����ψ���E`�,j�����Q�f۳�A�E��2��M�-��ᕿ�H�~��LH���C����ȉ��StF�Dwm�uL]�F����� \��F/������F�*NW�7n�+�g#�?��V��S�;���d�V�#��i֩̈EgӼ�ُK;m�����J�^�v7�E{W�kyX$܋��o��b��p��l�rY$�a�8X��XX1e{���}�i��O�W�5�'��98�)��K>"�'�@�k3A�97�'&[�V*GO��`�w�C�[u(Ǎt�������AJ��3 yt��Ο������X�V�~a	��7�f�jl"5/Z]�����+
�A����4̧�<Wܰ��� �X�*���)�*���M�MX�����2�e���oЍf��P4]�aa���z��^��]��Y�7it>bt��>��w�#�i�c�&��v���s���t�������%B�!�uq7"�����n3���D!�K$2��Z����Mu�pom�ݦ��ަ��8�#w����6;7��`����K�ڮ���>�J��W�-+��?�>R���;~���K
�j����h�"�\�{��Y?oz��n��V����
=ߛޓc�10��>ecf�Ɉ���k5!�O<i����G(�Ǚ9ᝍ�h��^e!�yשx�ꎜE���}�Y�Vi*q�~�"��4݆ ,��vWK���rGŎ���9?z�p
��WD��V� 蹨�Ax_�uj�E� ��~֙��q!�-bRk�Ɣ�,��5���c� ���sw^d��P��Y��V��=8&���FiɳSK����и��m�@#z������E����|��o ���p�4�f���%�o��z t�G�b�9s��vʔ#�r`�<b�(9b	JI��5K���Ab�ޜje��z�{#���l�)n�{R��v�4���[S@р�0�iU����8W���6�O�ʇ �N��ob-b�o� J�x*LB�G31��>�ET/�ƞ�D~����&�B��d�MN�;���?V-�ZP�)�1k ��d"ﾄɀ�3���"4�$�M#e��Z�ib����@��q�|5q4,�p���;{���㓑��
�[���1���͓rEM�����nb��:-µy��,7�݂# '��MMAj�j!��x���@>����G	���P��X���柢OP����X@,�-���=rn�c��	:�S��~�D6��)0gCI���yHHx���'����e��Z�%�4�9�B�xN!���3\���&�Ot�{��������'�Ӧk�vn�ܡ;W�ѐ1*�"g!�Q\=͏шD��*��������Di�%L@V��<dH,�h�t�&0����Lʣ�AN���&�Ė-)z��\����6�-^s�BS�ҥd��"�!�Z(��'�Rd�R����Om[�~BX����L��nQ3U���堉�?+^�
�]ŭX���E����V�6�[�\�g��5ܫ����G)ߧa�� L��i��t��&��	݋'���65~����+T?��!/4>8�e��rf�'_����e8�(�
tP��_��7��.L�V�W�;K}�N���ʩT�Db���Ӭ�W� ((|
g"�hC1�ɕllh�V|��ck���Y������`%�D�|�ǰE���o_? YZ�F�xƖ �Gm}E���!�$:��������>�����J�Q��x����0��\�N6�����j�΄a�J2V1Y��j����?�y��ʐ��s��
����L\�����H1���~�BNѰ&��4���M��b�굯zʰ8êR&�5��uN���9Zw����O{��ĲCi�$۰?��lK m���mݛ�h�(r+��g1�m��'�M%�R�?���6<�^?H�W� �I��z���~S���2��ɴY�q���#��7?�$Ԇ��NH��e���������픓ɻ
]8Ǻ]cs�/��X�N�G���W��j���xB#�^������뤫��'!qnG���z0�ˊ���W��}ǵLNIk���nY�>�Ȫ���� V&���Z��������q1�8~:�`{�M�� .d��^ �tA>A���u���-8� �x���L�v�f��{�!(|>tWY�}���D&a�ě����I�Wf�M,wC�$v���x��`��2�v��c+jG��e��J��Y�H��S�S����⟥Hatkt�V&	J^�̗���6A$�o}�<��|���T�F�đ���G�0CC���O���m4��_���%��w���;V9�`�%��p����?@(��A�Չ�8��>���s:�ˤ޽��={Y�����DQn��Q�wnr��	���wH����{J4���z�!}�/����~"���<�@{>� ����B0eq ��\]���Q������wcA{Z�0�8r튄���[#ǿ@�ȄLU:����5hh�s{�ĸ�A�2��GT?��T��P�澞�:��֦b�����A`����n�\�٠>5�ѩ��"���ڢ�g�G��}������~Ig��1����`��*CK�4��
M���^��!��\��7�}�oAw�b`IM� K�O��`57+&�q�t�g�+���s[��D	��&�����Ʀq]���	��lٽg.}����F\�	�R��pA�=�`�?�����P�y�^5?�ZD��c㇜(L=Ma�E���(�#�|�A�ڷt���Rn�\Z.;I7�d��f]Ɲ�o?���:��>�C�������$�R�u�q�G�w�^�j��_#RM�.,�׽:tXi1��y��B�<�n.9C��u$fhb�N����V�F�s���,S�U^�."m��Ӧ� ��+��E�Vn�R��%��zF�Ǵ���)>Ւ6�e��WpKgz�:�|�B�ѵ�'�[�]��E0qA+#u�|(��!�c�1h#Di��&����7Nx!�P�+kwϟ,3��
�V�/�G?0o�%0]]��i  ,P|���9�%�ƻ�9H��[27ۚY9��!��4�����:EHyށ�
�9;�ݙ�B>�+��{�Tm탦6r��w@������n�I{�<��>6W� Hb���j��p�s�@b�z�"цii9eo���j��|K�$>))�'�t�
�#�q�6�0S�y=.i�� ��r!՝٪�g�%h�M���bGGx!�rOj�2ög�?�Ee�Lv��*�La�n^��b/1H�5\a�'�a�@o�ct���3�3���T��d�x�/��2;�%e�fJ�-=_�oz G?�ρ_��c=���٫j�����on_~�������#h�b����K{�*����W����YѠ���͜=��q�^������-Ex��Mg屓�� �d�#�B�ӈH�uM/^rȶ�+� �R�L�Zv���0[�����P�60�����^f~+a��#!"�o^�9L��5�hG&(S��Ұ�6��ۣ�f�5j�Q�+̧c�6��@4Ё�N��hw<�[�Sk�,>ni��v0������������0R/%��"E"�X@�~7�R���U{�x�����C����D�X�fa�$):z3��U�i��w�P�^x�����\�E4�)h[�]
.�����A)��I�[&�}wf��n��8ƪb����u�(<
�fFG�^\{%�����[)��ij�e�1�{�"ƥ5.���~*�u�/ޥC*"����#��;��$_�5>֋��N�6��|�*2�c��/j#�LU.���ՍԈ�Ӽ v��8���e�-!�Z��\=�@5ή��B���f��`���[���VRD�g�OV����aQ4T� ��ZF�W�R�)9E��u����_���?��IH5���:�@-�nܹ�˞Z��h� ��㈺}�Z+��CG�V�����y��M��i:_3"��b�F����D`p�z�f��?=��J;����w��.�$�������L�j��(��k��R��
dO�iptG��hKi�����B��e �p����
��ذ��m8��U�_BS.�:�L��G��*���.���f��f"Q��v~�����p.gꭞ�|�0*��ɻ"����O~�:х\?��פX*q��cJP�Z/��!�n[��IPY<���|n��b�~��<v�(��䤂�}�s� �ڲ���p���D�C$��-%�,y ��Yɦ?�	we�^�q�����Z��#����pK��F` ��� V٨su��~����H��̴Ew�o�wbY�
��.[����\����*/�mߘ�#�*մ����]'z���Ζ�ھ�On��[L<�w��I}�kc��<���
�H��g觏��8�ӯMBf�}��?�3�euY������������P��\[k� �^$;����=]�f��U�U�����~��ç�'"��Ve:b��gw�>p��E��q���Qp�l���UU�vۧ��!��/�-l݅{	~`��O�� ��
�)v,g:�S���6�<���#QT�g�]NX��cc:�(��K 	����vg��Oª�KB]�`p�J�~���A<�eO���������5����i�i^�$��,�t>'Tuj�n�4�'����,�#v�
�>k��`���[<�acv>z~jZ�h�k<[�X ���B�9�֛X��+��̆�|�+]f�)���O���-���^ �n,�3RGe�SF���s�[�Ƌ��F�h�I����B� ��^#��1��]�J�f����$�%]*�q��P��)8]���|^����2d�cq:]�kn
N`�ù�9o,��B�ͩ�B0K^�J�9%�}w�JQ�
�ɐ���m�������	u�{XCA�D0���u|��Ʌ;�s�>(5�!Zx����#U�ј��Sg��/�\ST`D��~��y��0�An}���>��˛�,~u1uɒ�D� Z�'�ʲ4�2A�=__�8&�@E8��`U69�~��:탷ݖ�<���}%*J�l 0���f��?9�[�W
�(�#a��Sl&�c�C%�í�t�Q��a��b�:��$U~���;C:XpM��QڰL�oY�"���&�-��h2���XC4y� e�w����J�N$��0Z
$r�LIOK�j��N��	T�����	�7! ?��\o�獄��5#��9��5͍N����l,���Y���222`M���Xi?���J���F����6�۠�yKx����x�� �LX&$z�����b|\:���T񧇙_f�J�6���b��ȩx�۸�����G||����-M�=�ڤ��D����O3�R6�<��!����t��$��/�{��XCM����U+xV	v C6M`�@?�^>�8$�3ς�N�E��sy�0�_,Q�7�U���<�K2	9��e� PP��r�M�x A�p���4H�)�ƃY_�6��H1�ׅ��;�&:I{UQ2k�O%�k���I
q�x�O�2���FNM!+��۱<��a?���V���=B"���?d���7�8�	�ɌW�1ς��|#>e�7��d�%�$�Z�a{R����ײ��68d��f���/6�mU����4 �:�!�,ղ��2�n��
�7\4A�����e���-�������Pj�����J�q�$�y@�l���n�RAh����#��dLB"�.7T��J���_�PJ�B�T;� <�y�j��z�g\p�����%@��=|�CK�y	��=���+,YI�Vk���dM�%{�����Q -4h̋������h~"1�Al1D�����)�F�a�h��\�i�\�Cp,jG�����߷g��Lo!��*�����ȩm.EG�fgA��ܳ^���?'B��_(0�!R��x��v��o�m+��輳I2�(�뎒��.��g���s#�+04��L�2�XAD̜y�K��:��Ԯ!*Y̦hJ."���� �b��X�Bp�~l#~ʒ��2�2$�,��INx�p�r!|���=��#=و���M�!%�o��E��ч�Ba:nF���J�A����*�>��\+��gR�p�S>q��UǮ�mDfնN�����u�{Ld����7�� W=���7�k�X�ox���¶�����r�D3��m3�nRLm�_��ɀ���~���x�������j�n<������Ӫ���c2����m���ΌNS��ns/�D?U�%�^��i~ L��ľ�/�㱟Y���T y��l�c$F�o����y�*�<5qK!{�G�o`a鉵�AT�9g��>=B�o~@hwy�5j<]rq�G9I7F�5 	9�MYK�Ӹ�=���O�W���j�;���F�)��^�94��NŇ(Y&�k���M��L�66�a��u(m��^���s2F����yl�֣�7�,�2���o׀T���֧(�M��q���3͎��ڼR�x��^J]��ML�bB���q�s��N.���5���w��;���B����
�Db�GD��.uo��8�6�k��֫C�#���z���f�<
m���������P_���g�Y|3��Pd�)�D:{
A�\�����ke�&tX���lך��8kU+0u�S����)��p���Cʆ�G��Y����(��Un]J�؁�[���KÖa3��uq-��y{���m���R�@�c�ނ��`�j�e>!�c�x��[����Ӥ�'�7��Cf��"����6�G���n���y�x�>�9�r��V
5��qk� ^H��b�ԟF�?�o����3�������R	4G"�I=/V��8�45��y{�ڸ������Y���<%ݯ�#��&�&�~]aPb���N31�^�^���[��*��4����8�|8Gjl�5���Y4�Ή��7���[���İl~��п��i���YӇ���jw�ɘ��� �/ܤ��<�r� Ѓ1裶� 咣��p���n�EJ*�Awن,2�ȹ�����s<�nN	%c�s	�#�����m�Zr�q���=a&�dCgI� �k������@'K#����p#;.��� �_ΒD ld��гG������۾ܓ�����Qꔼ��Lp�^u�;�,L���]�W��J"��a�42�����e6}T��k��pj��`�>��X�K�g��H�~����x����miFw�:k��рjه�"d5� bڐ�v������&�b�=�Z�O�k��S���Q��s��,iȹ���qk5Œ��&C�#�=�.�w0J�lU�H���>�r�R`rv�J�~��h � /��ıZXY�H�-o��m��
�(�DX=3�s��B���fW
�8J�Mu�-��D2]0.��$$�܏ŀS��`P�%7�V0Wu�+�)A�T|�guO��m9��]]��>)�ݳg��|��%�Oj���&�'�q��=�X���\6��E��%�	��;�"eC\n�C$��8�m����\��J�|�y�a�A�����eC�O1~*r�V��ˋ��r{�}{q|,<�,֛�QE�M\s}�Bxi��mY����-i;�x�q%�s�\8����u����]Ly8^���hȽ��y\B`x17�?���y��Y+&s� ����&�RS�M �i��H�{�8).�����Kʓ��8��2c�L��
w�h���E]�8�~�B�0XUr�Wlf5�K΅WO�!�)%�>f�����uq׿i��7�*����,�O���N��2��+�CyQ)�#3����������W�E�[����<m�2��j<J<i� 
�c��F�o
���|#Xa�9�U�ZqI̅h���ojom0#�^� �Q��Ɩ��gA~Xτ���:����Sퟒ��6�Ht��9�_mI��~k@"�U	5�F�[@]m�~�*l�෧��$�]��ZW*b#��y�%Rn�I��}�r��P8��"1s�*س߽�Z�D�ǿGy����N����B�J�"��N��p
�&|�\��o����xԺ;��=���\F�*J��E���Q_�]r�v�.�[�i�`�}�̶�A��ol�!<⾕W^�6�f������M�"��d*)(�p����Y���AVȦ���]�9_��s@�qx뷇ٲ���!B�����R�u�TL�q���Y��`(�n�A9����-ܘ3�QǛ[I�|�F���t����~<�(XK*)��N<sرzU�;2�WCAE�Λە��UZ5�@�[�8�D�k��j~��\1��1�E	�Mw�m�#r ��0�7���;g1��e��[y�\��m�*�ZQǸF���h�&#.�R�͑�"=�,ڗ5%��������&�1wM7v����\_�Ɠd֞L������!~�!�h�I�UЋ�qȿC��">�!8jLY�	:���V&1Ay.`��ڴP����@^~�{6Zdy	�I���y0�3��fyT�]��WtY6��Ɨ\Q��_U�D���=!l��������9r%H!'Ӊ�h9�q�ҼmЯ<H���0n�US��: G������\�w�K�TLB��S`ic}j������& ��t��@�"͝\��>j�{��\���T�}�Q��k���B�3��b~h����@����Է<���Wʈ�fض�w�:B��&�#��-m_��"l7�@�U����ȴ�h��OnIh��P������j��y��[��':���Gq�@\�����)�-���>}X(>H��V�u�ul�h��{۞H��=�ҳ�e��Z����RX��ܐj��I�o��c�?2W�{���R��ŀ�/���}�F�����<p�ʺ�������&�ނ;@�j����U�Ч��򄙀ł^�
>�#7����>5��!`'B<fF�)��P�פ�8ń�\K1���fg���σ{�������!��r�C��jġ�NC�}�6��}��QJ�����.'�f� ]�/MCŇ�l����Eꀿ�C���%'��=��Z�H�
���-&�)�σL�Oag��I�>(Sm��m��P�W%Ye��ri�ɝ�Ӫ;�%���j�C���Y��<�A�
�~�G������&�R..����!�6�)LnزG��V�~��+Π�sV�_��F�j�������.���Q�up��RZ@�*;�{�e@Me
4I� ���M Z�2�)��z�`���E��k�ǿv ��كjh��[V� Q#��Ǹ����IR���5�O�$a���%Pdy��O�'RK+V��OVH>m
��o�_�溯���a��[�y�/ԕ\8�쪼�����e���w�?�!PXM-L ��,����	|#������B������E�똵�ח��$�E����S� X`|�7�Lr;ٵ|��I!WJv�n��U���uLl�0, fv�*��?MD`
$ �B�s����c���➣�����V��8��2r��n�5&��#������{�}�n� ���{H��r7cٱ#J�c��&O� ��Ă%�h��3?�>`WSdۧ�*�5���+�Q7��2D�'ٮo�P����fn�����P�]� ��]0��@�	D������L��Tc~w��~؍,!�CZ������y*�2,&��B�ɁW�.����s�O�C�bm�~�U[��'V}�͘#�r�̜)�I!��k2�t��Q� ��AsM��A|&㭒d;��Ĵ4�����a�ؚ�s��x����V�]�~~�5/�LYd�H��4��'$v js�p���^L�A���C�;�ӻ|E�p�%�<���c���P��� cW��=����\ڍ��x��a��3��а_k�����ݣ3T6dZ��۪���j�;߄�����ycg�x�,�re��Y��/g3�ß��
O2�w�M��P��gW�F�O�(3v1��I�p8��ӫ'����ɪЛ�<��~EP{��ň���V���BQ�Ҕ�@$����į0~�8e�h���.�tc`�7<9�R�/��&鬳���0��#ɐ(e�,Q��0��^+���=�(�������vIe2t��FR�[CM��,G��,0���7}S�R,e������;���b�����]������<�o�@�__�1Ҡ�<�������'�F#v$�Z���lU�2�fng�+�ۑ��r���1����论&�f�Մ*«:�^~'��w-��bd�����2D��5\=r�s��iT�#;ߕς0�p\�l��K�gI<�P�O�b�pD.�&���i��I5X_��$ �E�������Ab��L��G95x]H���q�+NV%~8SC^�S�.�+� :��*�����3�5'��&7�~���5)�e�F0��H�|���sP������ 6���j��:d��_fc!#5݈ '��D4�������˿�?�X|Ź��A$�E��7�Q��r#@NR!�#��I�2!|��u��|��F:9���#���#u�,����=���G�Ըcq���L��Q0 �W����Xڊ��`e�
Lֱ��nP��l^���<+�+�2�s�۩��V���S��悮s�{�~�T���;n93�x]�xê����̑A�'�}��\��P�_2[Ts� }�LLV|�3�P�%/��f��A�U�&����8�4q?ӽ&PtF��}�)�XO.���c#�Q�ӳ�F���6��S#ȱr��b�gK@2g�#`��ǥzx|��_���?��SB�M��u���Vا�����ۿ�\�G⟼�� P&W��n m/H���OX��]k��%l,X���
���R#)$�Hue'A��˯�5�AB	 �6�F��� �֓' ]�a�o���}�v��n���7�k��"~�/��~(N-��\��`l+���}���$��_s����J� y��S/$ԻDwf�v=-t�^"C�I�,_�c�N�â��&�L=��M�FB�Pv��-�<e^�H'XD�a_���i��$�0����@#�/�����n���'+t�?{�h%�<-O�e�}g�sw �b�$%ơE�����v�f�f/r�]nE���ޟ�,`�CZ�r5� �LEY5�aLH}	0�J4�@��(k�_�~;�&��E���N��ΗK�s70��ˊu�Ԥo��8�4cqX~	߇��sT��78�b�����X"�!��1��}�����m{ �h|���w�������>K���7W��OT�ӑ���S���Y�:4����iEw �ǈiS;�sV��K�䶻AG�#��Z���e�������Pf��k��>?mM�`GC��&l8���%�mAQ�j��N�����܁
�&E@�<�����5h����O�^���R+ x+�/Ƚ���3p_R���+�R�,D�����pSa8��D�K��(�x��5�ya�ک ȘXg�gS��:\��?,a�Q�Aj'�;9g0
���u�=����+�1�z�"��!�ŭ�X��2]J�tU�����GF�X(?��A���4�y,E���SeV�~[8��������С��1+�	=-�5���o�d�Cf�c��J�tų�_f�&��m���u�LTw��Lۙ�t��I���� <�I�`_2w�����/�-�0�pV����z���i`&�)�#):�oY�$�6�Z[)-�%ee2�b����l�>�C��eӾ&�&Q��t�}P(���_�4��~��h��~w�NK�3�?�`��v�\W�[��3�B$șҧ�ȑ�Me[��9�9op{h�ߐ����NzE�ß�.O��͇�n�wҹF�;���@����3o�!�����g
U�ڲ�H���,(�ch	�d��� ���~ވ�Ʈ�i��8OL�{��ߝp>�4[8$�_DU�:p�B�X=
ILl��C�2a����e�����GZd�G?-�ᳩB*R�'U�f�r���X��zоu����\����w-��⃻�K�ʮ)�&8��5ю����ѥO��Շm%���a� ��w ���~�"���)������wGm@@Z���º
T,$xȏ���?�_ӛ����(�H�0�X*",_H�!׊���;���������v-r�7��.{��V*&8�aG��CQ����ÓjH:^��oV�C��_m)�������b���Ç�ˈ��F���}u	��zI�cbcVIH���A �����f�!V���G�pDE1O�u�T�|*髰b�i"��-)�}���G�i���ee�o��$b�-�#~"l=H�42���W��f���"݀-��v��D6����04�����U|i�eٵ<�L�t+��Z����?:q���
'�p�CA2�{�W����at�[!�s>�W�Ә��}u���G�x�d���Ѯ��� GZ�5�e�uzW��S2d�U�^E����2��c��e���Ƭ�٥M+q�;j�%�<0(,�x���T ��}$�V� �ve���6������(�_E��j��S0uʥ�S3��X�h�S�T=g�|��L�[bOϡ@x�q�q��f���<�_Jխ��"���1ּۥ�?��,6�S �Y2���|H���)����(���2�v2�nG�)�{�I�On��դ�2��f{�u�|��<�h��4iU����1��hM���&���~�e*+;P�9���,mG���s\[�;=��Zo�����ӿq��������>��B;��(���+��e{}�+��_2ThU*��7��/h���X�|��c�:a1�hmt%�҄O}�Z��K�0*��!���|�Kb>�/8�c;�T	��kh�&\Sv��������)��K�8=Ur�V��K<Ӏ���O)"U��d��k�M> �����9+�	��:�	��S-�:�7����a�����^r65\R*<��՘�|�R%4C���:����y��W��"k�b�kJ�30=���-I��G�b�~�H�\�p�o�F\G��*�B3�K���܀ٰ=���G~��y�,�5����4�u}I�M�(&��ze�T|�E�J����u�m)Rp��?w�M�`�t��
�&��%ć��6E�^T�d��K�
��[n�i6;���ɿ��nc*��8:sx�X��dU��j�֣f /������V��)��o�%��l2�v�qT0�.n���B���T�Jn�p^���p'6o�S�t���������������>
����I�rN�;Ĥ�<� l�h"`$-ڐ?�&Ռ���e8Y��Uyf�'��dV����ef.� ��@�.�,)s�eIl��Z��(OUd\6V.�ԹN���;���]K����Iױ����� �x�9�]��-\�}@�NL���1�����5ڹ!��d�z�M�.��Ř��w?&"J�τ��][������x�P�L���9r���E��"�G0�W�([B�ak􉰴�+�&v�=�;R��Ȑ���CpZJ��I�s&g��5௩\B��*%�ۼ�c]����ꆥ�Gы 0F��,8�@��M���&���}�uZV[u�lB�܁���Ӓ�� tH0�G&�q��POCVD��"�Ԗ�j����$�?gHpz���B`�cF}��/9|s���I�,h�-CN�?�r  ��!��d$n�$p<BYQ;j���bܢ�9��E0��G��/Ah�k�i='�Մ����˫W>J��=�UY�I>����9���_��
�Xc0����~IؤB��} ҹ��� ~W�j��U[��S����9�o*���9��^E�_ij'>|3��y�%�.~il��e5�J(����]��) ��(����^��}���w	���ڧ���.Dz��}y0)�U5́\�Kay�t��c�gA��'�H�3������_�d���^h����6���朶)8X~0:P=~LZ�֜��cq9����gSIUڲ%�5��{�
�4d�\�>��+�z�l	�L9�"Z*�.�?˴	�G ޸���O
�a$~i�
�˲�����{�#X��u"���P��H��8�A�m��/�6�����c�e.�����5d2�m*��p^�_�ij/�A�Lzd!��|9�e1�����e�uwҹ�S�p{�s�����<����ȷJ�ߑdYy�1
�v�e���jh�%t7&4eƂd�u�@��J��(��#�_�>����Y��m��Q�-�0�.��E�'������=��8׃�$�2�eCr��C-� ϩ~�d}�f!��i�L���r=�Zo��AJ�v:��!==�6m}��YQ[��ν_��k�r ��޼��t�������H�R�/��{�z!4��Xq�?!<<x�a��Z)x��T�h�8�?����1��>b��oص���*f��R_X�0�����Ɗ���Tw��`�a��̜%uU�UPƖ+�dk���a;<��5[��RS��PV��'��O_|V�S!_�#�nVQfK2Y`���t��-S���d���q' @׮rzPw��U
�g�Wz��T�g���l`/�DJۅ�'Z����:JL%��}���&P�]�)���y{��;S�f���w�������Lme��X���Eҹ�Ĥ��dQ~�%h;Ð��3:�/�h������CQ��w+�P'i	��������7�� ��]�q�?���,�[[;%jca�U���h��ɛ��
��������^F���D���`Wq��WiRďi#��(������K[��$G�G"A��b�֯�eD� Wq�]���T�%��d���1`{j� .�w�%թni=Z~3�Z�q+��Qr�<�k��b�����;Ŭ0)�bp&�ڮe_+V�K7�6{C��c5~�l�.���4t�ڍ�(@�8B��7��?lq��	T���ۋ�b���V�'��A��Q�RU�c�dy/���x@��������3�����T����^J��	>��pdU�9R!TY ��)��7�H�Œ!�_�D�G+y�Q*<�.5���\��VÊ��M���4���Ӹ�'j��G��0�څ��r��u�x<�^�w�؜��6~8sђ��
�9�2j���7%�ऋ�#�A�+z[9��l	pe�ZTM��5l��Km�2l�N��8�H��*%s��3h�������a=�ң�����	/B�%��tI����}'��,�����ǲ=�s>�)W�z������"0�|T�D�ܼ\T��p�S�_�]l��3;=�VM�i��7?�]9�C�B�zH���;�@��O��
G\��E��0�-�~��\Q�s��w�@]��Ƞ�j�)"fȮ��R��)�kS�yj'�� ��ޗ�Ƅxj�N�A�����3��3�3)ʡ0�s.ă?V�������F�m���u�9wR\K	���I��u\oL�W�p /���d�
�B�GX3§Z�1+� ��"�	0h��x�r�(�&��w��+�Ӆ�X���+J��}c��~��)[�i�f���#�������#�/�z��Lf 59���[�g��XJU1R:Sމ$¢;>9JꫣV��TmzP����l~:d.�Yдo~!f��$6Ig�a�n��
���Q���\'Ώs���k(�?6�Y�V���Ч�HC�]�9�V���4�`��n���Aw����
�������@Ф�Ż�T����#��.�IW���&m��0i����-a�����:�ޗ�J��xvI�39<�X��r~!S����V|�sh��|Ѷ"��7���e�[uS�	j���el3��V9�}d>���K㎸�JBL���y3��;��j.~��Fe��Sy�����"�(�1�6��&w���Y�ƓPц�I�'y=0����Q��~̗�YUP����}���#��B������a��|v�0ܢ����$�E��+���x��2kٲ�NXNэ��rV�g��(I3:��b��\��}3n�FgI}P�R�2�f��01B�0�S��)󮰃���G��RI<ϲa>���5����2l���hp\�|����~�CȀ{o���c3�n����	��T5N���W;�$b)�q��E�+���OG��˜�r�oy�	l�����Wd��j盻Ev��S���jq3�R���b7��ǹY�%CZ��P�e`���O5�I)��@�U�{�W���2]�
η�0 +��*������"}�3{��>��0 ��5|B�^x�\	�q��C��fH����B��G�l�F���5mB�:ZTW���z{F5*�_U�=w��i8���E��kP�.�}�t��rm;��[�~��
����z}��S;O'��?�����ez��nWFȹ�ߙ����M�R���<�;�NԿ�ڧ��xׄ�S?z�a%- I����n�1�n>�P왓^��l��Ӆ�ȭȞf;�R�!��xc���0� �\��k�k��s�f��ȅX		�:[\�UCK�dhhX�܏e��V��{�����v�q��n\-��h��n�|=)��X�ڮH�5��$��Фž��G�s����OG!���r����ʔ�C����Gc$�70Ǳe���L���OQ����<,��"u���u������t^|6i|ک�}���Z8 ����M���#o�e;��1�F�u��F�l�	�X�Q���Z)�*��<%�i�خ�h<��s�x8Y҃eɰ|[��)��dD6(1�(�k/���[ۆ(���������6�F�����\�˒y���4��+/a�fE_$ ^5�vF���b,�/`W5��C�t�rrt�8����7��8&�`	��**A��E��Q�g�s��MpdR؇~8s��G�����ߣ���L���� �e4��[��3��©�㩈$b�x��eJ�Q����Ɛ��Ψ�mmÌ�$9�{����=�%�^u
*Ĝ&ji��!^k���42$s}�����ta����n�Ow���-<�*&���rz�>K/�tTT�{?k���Y�0��b@�r�\��Q�5>���iB�oy\/boVF�.U~��Ʋ&R�n����fV0�b��I����Q8ģ������s�˯���������{���)�t��@�fq�0�R�	$��ӝ���CRW�N:�ٙ�|��Gqyf��Q�[c��M�CKY���:���~�# ���)����5k��t�E�|�.���r���ۋ@�����e�d钟��,��V-�lߛ
)�l0S��y�R?tf]I�9��t.�����Z`��?��0����t�"��Ne]��.X�)z�6����YfW�a#]Q���Ja���fvD�� 1ϱ������3A9��n��INB�%�cA4:c���_8-��Շ��<Ä�a�5����1�q݇vfU�N_���Kj��'�6�iQ�3q}����xw�$ѿ��TT�QQ�|'�(mGM�Q��vǢ��4g����t�+֝������%�ש���O��'��5�B5��_�x�\��v�@�,��~ȿ�'��p�pT�>�U��8
����X��`��Os�릣�Jn��|Yd
;|�%ys�U�b#�vB	Q�_��9��V��T��m�5�ŵ�{q3�1��C|�u)e=9�:+��F�ss�t�#��y@�f��>Id��h-�ӑ�0_���q�,�%f�t X�||��A6hcc���Ji��I.*�='/�~�W)\`�/�;���F�pm���)�.h�Q�X=�!��%�G�$y�lH$e6PܙJ��`ͳtb�:~y�/r��Nӗ��g�SP�!9ы;R7�x#3=J:=�)�6᝸G��Gsk-7<	^�����'�Khk' 9�<�H�CP.k[�!^v2��������u@�� �)*�Ѡ��6�X�`!D�%'�~�W��>������n���tS�e��L�!�U!V�W�F����i���&Im�խU'f�Ţn�J�Ř{p=K�l�n��W^E:����ZG�Q�//l#�Z��C.X�g@d�?o#Nܲ�a7�-��������-z����ě�l����UŢWOI���Ν�2���m%9�����eH���ڐu"��<}Vw����La�Q��2ٺ��s�Ϗʌg�hi���*x�`��V��\��0�Sk7������	�5��ܸ�,�".�|?A�1>�ҷC�*D��Mr�\��{�u7�0�s�I)��ǔY����{X��?� b+�5A'�dfb�{"�D w,���Ml�۔k�(s�/�]�w��#�2�����k���C}��Qr�n%iz��k�e�G�%��-�󺟑�!�	#
lk�J���.�w����ܤ���RT�'�D2�t� �.����ێ�d�h�f��}�k;��C�	��%x��'���i�9bY@��Km#��]PT�s�s`1`a:�3pBĪU�����貋�fe~#�T~Y��ޮ��ż{�A�xܑj$���s��m]��E�Bl�3��}�W��Q������A/Ve�u��i+o�&�>���판�o��v5�����h�w����R�=��EkЗ�#L�����(��]��u0��54�j�YN�k)ϲL��<�FN��j�s&0B �G���m�t2b�H��"Y��oY ����Hڈs�V�.\����a�n�X8&�3��4;,���!E��}Ly��[���gp�	%3$�b\��~���qnp�|��
Y8���+�F�j?�49V�������C�Hxs���(�6v���k�?�(F��&����^v������$b_�:��։��5��*.\�^X@�t���DB#�薥+R�h��3��۞l@.��{��&��Y���&���+z��8Iw�"k�����0��J%qy��q�7�' c�y,�K�!�-�ƭ�ӀƆ ��V�d�F��Ft`�74.�&�MqٮY̑��� ����}�C��a(��`�y����ԁ��E{G��1m�b]��mٶ�auY�iN� ������z[�_Xf>+��QK����a�Q�=P�	$��f.�H��t* ��<�8yr���O3 �x��Xۓr�՛-яN�N�S�.U%c���3��f�#|�7�����A����1��{�pW%��G�/��0?rY�ϛ{_����t�4��QKi6�]QCc�_��=���&�(�EܰI��|㵄}�����X���Rx\~Z|�}�N�>V��$��7��h��Az"�-��l}�H9�P�5�1��Q�Y\ /L���6 �ǲ�}P�kv�g(�(J�!}�Am�����*��=r���r�<�E��x��^��*D�ѱ�=%��9/�W1E"l&��*�:>�'f_v�BQ.�� �!�4!dJ�i��eY,�η�����	�ii���h�q�51����[djC:�\T��%�7s1��;�5M(i���Y�U/��6��j��K�!C0!p��q?��ݎ��|rr�>�Ӎ�bV2Ѭ{�N�z	��z�h-��/h�J�&� i�k��� ��u~]Y�m����I�������:IG0� nuvɹ1@v��1�>4��&P�v,����\%^dv U�Z(-�X�њ2�^�����!H́8�hM��Ӻ�,�#h�oG�Q\�:9���`uSVֶ@|g��J�����tT{����H�:����e��Ӛt�j�y��2`�appW$rC�K�9��:��̦w�O�MLZ�s������`�V����OJ�!��ƀL�]T�߬��e)�~7ғ׫+\���-�(܁�C��'�`w�=΄���"wħ'���'8�p��`bWq~��D�����)o��Xf1��*GD��l�k.��e��L�;�?)3��L�Ҭf�z͘%�>*)�� t�}�~z "�}�\B���xj�sJ�V�U�D�� �r*���D��O���C@%���(3{��/�O��䕃���U�ɏ����)��N�$��EgQ���g2�r��$m���{�vl�j��4xs+�l�;tv�{��GX�of���/����@YM%��x�9���!���3_�bj���a�@�q�D'�*���R�#���9t�V��b�tI���җ��Ø�6��]H�t�Jr��20�"X��*��ik�B��&�����ӊ>�JO�Y�H�e�u:* �`��;�(����PLu2	���
�ra	uo�N�2��%��)�lYl;		����c�g�{�D[��m�V��[wQDx�/��N��ni�M*�à_����p� M��;@]6��-`�6/mF���-p�˟zl��Z{����Xʙ�\�	�`2��I�P�&�(�5PP�y�P��w�7��yn.?s�
�<Z�|fV5��T���c��·_�"�9��эw�c�:��s �ޫ���5�����p�G�X�ǁ�>x���; ~"�Ja��ʆ�/<OPH��.�ow�O+���%v!��e����z�e��Vَ��f)F����������?�*�_�ێ��N#W0�Ɍ&7{���x*"��aP�	�ʷv��9?�e��N���$$��{�h��ij�tC��͌� �
�6W�S;��?v�6�4�^ÅN��J_�7�^�~�t��`܊M�=�(4y�OP��?���6���8�k� ����ag\�pg�mR�|.�jϖ_�mE��8��ǕU�*�K0��"��\���M�c��5R&��
�f)Y�5�	�.=|�UI��9��
W�@����͠���^0��*P��f�(�rs��4	"�%Ϥ#���J�����!�Ј�NF��1�7U���O7T���	���UW���alv%����B�w���� Ѥ��N�F?J]V�.ÖpgUJ���L
���]����FԙΎ�zU^���'C0�g>(:�d�e��Y#����;G�i�˪�;��9�Sd�AY�pҟsD��6�)�P�D�>�@�
���wy]2�O͉b���5���>�V��9��}iN���P�������t�y/�c�}�s�gjϛ��)��CuJa/�W!�?��pY�~e:'�4Ґ�g��yjIr l7>��t.q^�.�licѪ�Uz~4mv57��69KF0e��9���j,���XdN�^wr��f@���	`J+�E(��������"KVrĕ����:��Oӭ�4�N��|n`X�� k�nq�[$
}����E����Wո-�pR}���r���\C�u����A������ʾ��i�R�,�"P>g��<ߵ�����?��,E�/o�d�uW��Jf@�Ĥ�^�D�'D@���{�/ޖd�@�+�[*J!��`]o��UFvsU�Ӫ�GWn�����[s�lE.���K�s%.�p���@�����)0l�����t������5,��j3c�r�[
�Fћg���zFkC|�����n���-�wGyV��op2v"�3<#��4�-0�<�M��O�r���Xӊ����]�Rr���a_6�jA7�B�4,�
W��;�s��V�m4���'�ꮣt{��gG=ً�y��t��e:��C`���p�����F�CY���{�ν��q� �& Uj�z-������~�l����I�>ߍG�����#g���~������1(���2�e���D������=�*��H^�*8�rz߻5��غw���g�I����(��]��<$�����IS*J{�sC%�/��3�!��?�I� ��&Gm�n�QoI�i���u�hZy^+}؞5��ʚV��E?ᖳ?������������+������F�'�&Ç��UY��E��&�/����Z�Idr�3��PT�P���;�E.H�<Rq�?��+���?3\{I *����0wK�r%q��l-j�p����,���[@x�6H;n�q��X7w���O�����f��	�'�M�穔���ɝZ�`�|�CAT�W3s[����?+|#a�].ԏs��0OЖ���#eЋ½��tdX��XE�Z�S:�0HA�>������ _Q�F4��LzW�&����ܿ�`fr�D�N�7��3)���̨'���>rd�[��8t�;@_����oW�@VA�n����I�D׹} �� ��x�O���y�������L�b����.��7��VDe����&�O�^E[��\�T8x��[8z�M)�y�V���s������a"��	�ߖI��Z+J2����U��Zǆ5�ueOm�D1�}�	,
�Erfbj���/_
�E�R�85;2��b@�� �Q�:?y�{��H��,x'g�- �;�r\ѨC �8��E�\�g�d��Z��mC
�Z��8�;y��lf��D_�����h���-�i���<�'�1Z10�0�^b�HC�K�6�3��ۂ�'�M�� *���b��KC��g�N��86+�+� Ԣf�G +�E>+PA9t� T�%S(�'��*Q(.4@c��5��T!Q+�[���{�!5���J-"Ɨ�f�(� [C����B�ē�^���*�^М�(��(�Gi*�St�J@�
>�Ic�z�ׂi�y"iȻ�S=]�J1�[���$e���$�[zd,���E��=߼���A�&�8]��5=9�;��=� St���4[�����?�>&��Vߦ��S�!�d�bH=�GUp��m`' �ejȫW����]��� ����N�ŏ9ߴ�g�w����L��ϧAwٝ��c>!��f�������Yy<��BP�|���W7)�>�mLd�d!M�Q^=��J�����\�$���Z�
�͇xi���e��F�^K�֪��0
��Iy�C�Q���f��>��0�ޝ���29먇1�*c@��r�2X΀AT�J���I�l{�(1�!�����xT��W�d��� ٳ�ש���'�,o][��"a1Ĺp]ߵ8��}	(��� �wP��C/"���M���hPNNG��^شk��vҩ��PXI�ɇ�H��w�h�X�wJ����b����[}}IG#.�����v8#�YԺ�����1-[I��Bl��$U���L�3�)�y6�2�_��_���8&�Xn�5���ii�aҙ�	;h�h��E��'_f|��Y�+��!Cd' ���%T�f��yV:�UJL bE}J��R��{m7�8*�d}qi�MQO�_=��`�t���
`g�za<,垓v����`��nIX�O6.M��>Rq����]lP��P��1n��	}y�)y��/�ü����Wx��W"p_�'>�����3�2�O4T��V'*B��u[�f#��C�i��O�5��	E;�iNf���X���60sk�7XTB�3c�5B���Gg&���d@�Qbi�?�&��8�L�u�p��������w�pj��220=���@���O�`�`;g�<ڐc67�W��UHa.��p�#b��S�Zw�~B�AFq){�͈\fr�5T!������h��Yn ^	+(c r$�����Puc�A����i)���=�]�>�R�� ��w��?7_|��*+��4���dH��7�T�u� &��P�Ԁd�;<Bݏ�z��\�V�����/1���-�� �᭒�׀��S9J�>��g�\���@^��0H��jL� +��3E~'�8GG�q+�ʇ_T^[-je��=n!�Җ���W���*f~�&�Yqw���5s����̊;8���=5}!i�>V�]�%��Wz��gca�8�;?�Z�qkhD4����;m���B�4�����Y2����������Sȿ��q�nJ���a��^��6�l.[١��&���/p1Veia1o��ȇ�A帝���>_Z0�)im&7���Ġ	�L�P9x5�������G��Ys��+��0���Ȫ��K�,)#��dc���s�'��q�¸��Ib��E�Pc�II^�s;`nT���e"0W4D�ɫn�#m�-�O*8�S\����N
F�'��o
��½6���G���\:z^\ȯ���\�| ��~�q߃�9�S'��K�Cn�c䓥�h�~Pu���2/�����a���[�bt3\�g��9�����gY,'G�a r��L���H�ӹ�%H7���|,+���p����`��$��JS����~u��i�4�������D����W����I�nD#�v��S��a�JJH�g�w^��˫�z������ߚ����II�""��߄A_���e�׼UT�Z�Փ
O�aօ�*	"ћv11e7^�{�@2���M!:��--�7cT�E:��HZt���X���������߮�,b]j
��s�����̧��U�.��Ϥ?���|�1�.EРN�n�|�eH6��&��E�7!�)���
��[)ǀ�H��0F�JG�f�q�H�.8�Q$����Ӣ஽p�|F���	���݅�}�Z����O�	Ǣ��@$�)��	��#���㰵��IK�/5�!��qf`Otc���dhBÍ��YNP[ӎ�%�n	R|���N�.�\߭{n5�|1v�@�5��r`o��XsđK�����]	.�
f܇�`}��u�N�߻"��:Қi�9?N◠��
��zu����fF��ש��a�'�(t�����]������e'ã���<�0���D���apU3���2;�j׳�x������##�s�~ǋi��3<�L%rDe���1eWZ�`��H���3���E��1>W�]�`����&@����5���~���XZ����t*��Mlk�F�ϯ����XYu_�GM���p���H�P�|�Mn�	9�z���+wd�� ~�����b5c�ٖN� p'_p�Ƅ%'#�Gz�B�J|��M`Ƈ]�{�]�%��� <SX����N��T�qP�y�@P�K|}�}������a�j2Q=�28���nԔ @HP37�_y�������)4��Ē�<ci�Z�t�VTx��͝f�𤓳ш��d��������Y��.n�qc��Zg;�PQS��AXt���Oc�5kC�̿%��ՈYj-�6V�7J����e�,�D�����6BH���*�@����Wyl��TȉX�**�hCn7��qP�(����б����_�;L�9��?�o���I�ps`j6<������A?�>� �±e�  �"�QY��a�B�藚�����pcA�k���-M���|S���,U��S,�ڰ2CG�|H�`�˭;D:V�0��Zu$��ϵ��B�4�1����l_�����Ȓ�kw��sgzbU�$�o�eb8��R���+ ���d�"#��B<I�2�/'D�f�d���˥��n��f�`�Ԗx��N	wQJ��EK�My��i��ն����'��w`'vO5�ᱴ>}_dK�O1@��E��$�p�@�c�2[.ØeO ���Y9t���Tʏ"�A��PZ�X��/Hj�~�$��K�s��'nv} ������8�r,�v8�?l	]&�4Փ
 ��)J�z(�x ���8U��&��S�3���2mBB����U*��n���|u*A��gYo'�Q4��E^�f}�W�3���;[x���@>Ks��1)�x���ֱ����%� /��-�o`pVجm@�}U煈ML7���x��4�@�PH���Յķ�����>��UVIM�Q[dK���������V��@���[Tj�}2��p
gg/�Ƌ�ޖ���m���na$Nŀ*���OU���?25W
���%�q-4�86��u�ߧ��j`����pp���W��l88٬8�2�A0I�S�V���jp��#��S��E�E ���dw��	W�)�,�s�u2^��H�K����㲹���vH(Y#�^갑���OyI�q�H�Vu"�`�,o�5)������(i�ɋ�.a_Xe�-�M"�o���]u8��t|�z/��j��J�o��k��`��f ��g�Hޏ >�z'��"��6�m�t���Ħ�&4����XÊ#d����Gj�����s2R����NK�T��^���eU��{-�upQ<�*q۝i��R�8� �<�o�s=l�#C�� Q}��@�i�@��r�$@�/X���G�^֬���ẁ�����G�@���5�t��$=���]SӀ���e���Oq��i=�j�2�;�mۻ�U�u��?��]���p�#����¸~�p��(���z�U�0�5�5�p�N:vt�����6��r||_�9p*6Fe�Ȓf�?V�}��n*W�A�Ĝ�ԝ�cH�y��&�t�I�~�KQV����h$"s]vN�����Bs2oG~%cY�%p*��e�>J�q�;��������x���l��pc�x.��L]�[Z'�*�<�H�X�,}���*V��������>On3R�A�~gYE�x!�a�|&x@� 9ϴn]s51b@�*$�KK�[؃s��{ov�����/A�}*�H~�璚g�_q4e͵0��`���VtQ���W�����P�/~.��u7偬��)��l��Ƚ������� _b��,����96�`����Op91��y]ۻ�O̤���;D�d�9�{�*ZE6ˠ��:�H���8��������a�{~J��p���.`�^5���3�TgF�>�,}®Y�4T�]Kwĭ.��6E�?՝�u�FY8C��B(ǟy��7]���_���JM�0ðu�\a�|٢�q�J�oZbav��� �c@��[�����L��À�¸M\	:0T�;�Gڑ��2Nd��氰a�b��Â}jXJ�Cq7^�cCUk]\&�$.�Ű��w�C��nzi��3��̹^��*I��(S�˞Y�3�(�6�o�8�t�򞠎\f�e��b�RZ����<�.���͗��&��Y��m�Ѳw�s�,���a⮡��U��,/0�9�'!�ЅCL�����VH��`),D�](��!�$�M��@8i����߁ ǀ7�\v ��Y��"�3C�mQ4J瘃9x�5��Q�hw.��Ӭ��_*~[�����?:N�lq�� X%e :D�.�Ɉc�&��%�g�R)���Jj��ޟH-�USWٸq	T�]�%X���ߨ�#�$�-�cKtG�W��r�!Sj Gp�A6�&��n�����eo�*���Jp�/>�ךZ�7&2�r��k�cM�ьcu�|տx��9�Vy�N)+�xl��2��-<��&9�o�ִ]:~>W��oE�6q&R����C��U0���� ��[��̜^�ޮ���d��N�_/��z$�����)MQhv6z]]���*m�+%?"��qL�@���O�w���d����\~P9�A����aڀ��`̧n>[ȶ�*��^��U�	��iu���̶�;�I��sZ2�,Fc���I�F؉Fp�M�l�/�� p��4�n<U�m�#��Od�WYHm\}�ql�u���L�{�9�E�ӓ�ݰ>@���F]�)���q�H�)@�RZ�qd��s�uff����U=ARL�V�梺�t����C�ڜ��0���L<�������/�8c�i�����M˫�XF;N�|����R��6�.�燚����2�AW�����ä�}�����1�[X�?��h�4�/��l�>q�#4NN�1�#���߃�<ei�ˠCco)z��n���Ӿ� �p<1.��'��uCJps�a�ӓ�xT�-�Q���E�ѓ�;�ȋo6���S{4�������.T��Am66Wc��Ij,� 9�"@��g.�x��2N��0]�z�l:�fؾQB]��yC���UQM_�9�}������$Q0r�1^��j��`� C��&b�4T�n�_ћ������C|`����Q{�vϦ�F�qG��\`��%
(8�<@��B-��	�mj��" �X X��	��W���'�;�v:�S�����1Rn\�	ܞc/��iӿ������I4�_�%�b�����t���wf���$kY���$FlK*�\/aI�p��~�������9q����z���i�c�R�oaa�9W����
��l�	�����
R�{�����i��⊟~�16ΦN�;@RiDΆ�xlbO4$V�2��� ����0?�#��~'tMP����A��}��웛o3CX*���q�u��c�Ͻ@`%��W1��.Կ�A�(���紇,�w���r��ɑ{���CήS��%��J�|��d,��E+���[#d3��I��+TXz�]���Y'\�o��J��˽��y�*���
C~卶��ݨ��<������U�x�\ؠ�DC�֮��OR)2�>��`�YvZy�HR�nc���;�
�'�r#���S!�NE#�t���lP>G��,?���J���J�&e幅��2JˊV]�|,��6��v�3�hYЫcR/dR�/M6�G�`I�u��m5�UW�}O��!	�n\&,��	����W�5hhH��ꂑ��3�@�F�Ŋ�?��.9���لT�~�*���Pm�M�!�b��u�^輒SMv;V�pF��!�gq���ɓ q��I�e���Sc]��K�B��g�W�����+�b� u:��W�plVD�p�pz(L�Gb�LF5�"�";ц��̵�i~���Q�t
F^ލ\ױ-\���P�T�z2J:I%����m�U��Y�����?�U�|Q#I��D]�<uLwp"
X�CY�6�^6���;[�N�܆�1Ĺ�:�>�ѪU�Wfʗ.
��F\�"��"-���
�d;�8�y��˴ybI-_���.6`N��V3?�t�9�1�"�+@��T��Nq��|[vc�Z�p~���.zf;��ph�n�`�zr��E{�������W�ImXr��c�t���ƚ��f�����1]�lw"�)�q��Nj@x�]y逺�|���v�^�k2�����u�@��O��������f>B�Y�����;�5_*���26D�
�L�E4�"�+������'t��q�� &e��� ':1o���;M3���,����+��H�K���I�"߮���e�EH[��k�M������Zd�?2G�x͊.MS���K
25�)���@\�'Y��&ޱB
����*ycDP̶��yܧ�.�������co�#��l! *�|����T!������*���#�q ���nN�����	XNq:\3tR"�I-���X̩X�|�/��������X�{rQ���n����-�h�p�six�`4ߤ�Ko����[[�F覊p1�_k���#gU�H��D��p��?���҅/�;�����ﳼ�5�[��%�ؚ�]���a�(����$ϼ�_���I��Y�c�K�s�%��p?&@M<�kC��>�BH؊pQO�l��������]Hk|k�a����W�d�M�����&�
�My�ʲ���@�SM�#�P��T\=�0%���IBC�ň�γcq�k������/!��=��,������)�cq�:�u�L�91(�г;͘�X!RJG�����.WW�\���
�	ЮR�r���8�}W����D�H�0���u�K�MA��&{j��${��d����O^��L�a�w�HYDeyly�c��TT�HUY��)���>�KnX'�,L�[��ႽB�~{|��7���"��ʛ#��G�
�H���g"Â�J��Hq`�8�@���s]���e�|��p��p]F_��z"δ����]\�|���Rx���-� q�?�K�V���oY	6�ϡ�Z��`���)xyiA������=eX��*����a�e �V��'���LQ%e��j���Z��r܋�vn��ƮF�={�z�l���=����RI������I��b���_�C��V�\;�9�a,�6���wW�ő��)E5	�{5I@.�n�^Ym�>���|+~(��5�r�WZl���rGP�`#�,�����y�#o]����Vs gQ���LWO
�%d"�>"I%�JmfН
�7R}+�P 6}D�w����+�`�|h�6^y��#�d�3��0����cf�_a�.������c@n@"V0ʙ��y�zk�TR��gY>����o�tI'�|�.z�?m"�pω[$V���+�=.C���V�K��挪H��Ce<���Bz���N�2�O��28&h�DI�F����%V�8�d���<�1o��E�C�_��y'@����U�'8b�_U�P@(��?>�Q��"|��S	��-����rüj���' G���q<���"2����]q�^��=�5�,���La��Ƽ�g�,�=D掷z���tK����f��bj�ɷ�:mŃ���I����<��L���HoX�bi_�͍ן�eI�b�b�s���yv��Ip�yW�N�-�k��K�?���R��%���9_f�B�8y�o�",@�:]e<樎 (�)T���-@M;u)m�ƱDL1O#4���$���E��/
i�
��
�!dk=Y ���+�A(�^����g�Dr�/��T�;�ʫ Ik����`�����"@��⿞Jї:��ArLiQ��ؽ�����5Nya��V=l����]_�Qz���'��<�bwa��'��4�ϴa)ӗlx�� %<�����S�N. �<�DH�QSw�ϑ�oۈ�)���F%ɮr,o�(�f��e�5��m`+_�7q����$O�/�{-Ə�슣��sep��>ŸQ?��;�_��:�p���v�9�|guI�� ���l����>�Gj�%3`�&o�3�D�(.mM�h�l}<اI"��Z���<4��˞�����W�K���u������l�~�MJS��^���r�O�m��y��KadA�Mɉ���a ���D�2i�`��K���jf 5���R��k���Z-��u�{��������́���IJ�A.|����p�6D��q�J)�2>�Ov���Ī��Zz��K���.>�<�`���h-xw3�n��)���R`�PeZ�/)�Ax����\k2���c��N��
���M�wF|���j��[�?������a��/�/f:#�EB�2����-f�I��ń<�$U����ٽ��o�����#@�ݼ��녩�Mun�l������L�>XЄ9���<�Pv�W(����_�R��<wj�љ�ؔ�g��i�U�<�e�!̀M�2�S�Xظ�&��\�_�6��X�m���@Ǩ^�?a����Ҁ��~ׄ��+��K��i��2j�����(1����8R�G�Q����#�{z�1��u>\eּ�g�9��6�̾�~��'7Z�A#¬ C�vYL���c�/ׁ \ݩ�����A�p���?�s���xo�}�\^4/��J�W�=�B�!-��M��Uu���V࠿k~@T8>�v�</��;�!�six����gS��o�����_�=�WGԔ��8��Y�
^��b��Hq~&�ةy�P%���GG��<���ۉZ%����(K�*�������j������x�v����Wq��"d�6������ ��d9LY=Z�uV7Jb���Z��Ar�{�ѱB4��� �0���SoX��t��pS���8T�6�**2y��Ƃr���D.R0���,:�`D���j����=&Z�+�J).6��7@%f0G2��<r����	���W?�]M3�-����P8�M��R.g/KuW:��Qك����%� ��|ZB-9r!g�[i� =Z�Sfz�<�3�G�WSb���_ W�ۗS��/:�1�HbM>���;&~mmB^�e�qK����~�M7����� ��O�ҖzGF����oܗ�	g�����
�6q]�9Jb��'�x��H/� Y�u�h�h��H�I��H��>C�W�I[k�#�>w�>۵~�$�3<���!��G7_�=4�=�-Ѿ�U���(a�nnl)���ӞX jI�R���0w2��Ǝ�&#�����F�:-q�c&�o��ɼ
J���}{�m��/Ĕ�s��v�#��gH5�x�8��
𯾵h�1����k=66�NZ�~�d��`�F�&df�~�P��Ss�)u_s푾D>[C�Ucݨs��JZZ�a���ø�(�t� n��M�xu���c/|$]�"Jk����y�,����{�&D�s!���6R�q�d��t�K�.�P�q�Bvy��WL�Ԓ�EZ�GE���y���]���E%�w$�A�(�Ĺ�̶H3��b�Dv(n;�n3�u��jiA�՟�;�#��-њ�n�[}9�w� ���CG���� �F�2�+���#�~�,��߄Z����^4M��p0�,J��h�p�e����؉����8k���EA.k�L�y�L��)�u�~ܮ0;�cC"���U��
�lx��)]i��#zz����r].��ڇ��<���	�A1�*n7��
��,��Y;�E>�`P�c=E��6����H_.vi��
DqaU���~t��	��8���M�3S��C.w�����k�g1v-6��Q���-{���� ņO��B������1���ǥ����'�)��3�>C�z�@{go�'R]�p�o�*�U7�+�[��D�ڒ�ÜЈ�?���j���Wy0�Q*Bb�jq�`깤y7��A��yd��s�GŮ�y}�ׯBn0��l8|u#K���m'{�-��9x��I��M/���FtÇ2���\�щrdp��1K��A�865U�h�o?����pq_��?Ґ[􃢺,�SJ�jK�?b�Ro�t���. ��Xc^!%��=f� �*�8��\�l�n����axhln�R�4V��ѡ%r8�#[�%���������DTF�ˤ��:����9����ۻR�VVAv�sR88��J��M �S���E�'���K��"��(�C�4��Q��D0K�_>��"�ޤ3do��r�#[��Wc�*Nʄ+ڀ��)#�^SRl�����)�I���Ѫ���悱�pq�4Dy�0f�8	L��z��Ê�����p��V�):���A���n\�la&x��{!L��R�T:\��&3��1B�{Y�uOYM�xcL����(
Z�����s����C�P{w�?LX9���C|�%�s�u1��N2O�w�k���؋��!mEES}Yq�ϋ0�'t~��I��p������h���+.�-U]!%�_l�����j9B�O�O9�#�Үm]���������p#L�fg>5�f��J�y1��1��[�[_�}�\�4��M���|p�.�L�vdV�6���#N������!��{��xS�j��]�-�z���>_�d��V�����eG%�!�<�s�g���o�L��3�MO�fM�]gə��9¾��/|!�#�I+�6���K�|��S�I>�yC���+/8p�O!,�^	,�3�Mk7u�rB`�UW�ؠ��m�o��G*h'���VlP��O���B�ٿ��=�ڼ0^J�=>z�����&*h�ܾ��+J� K��j"�+��d�d?Sr�w
��K�D!�d�_���(�d>~6�bӳ66�D���^�k/(�|R��/a����o,��w��3w�k�z�SF�,sS��M��z�ͼ��3D��E@�q���)7�쫱�Uh����jR��"�Q��(T��Ȝ��@�~�IR�ʀ���[*Q%�ek.����d��7Tw��PR�%Ӌ�o�Ag�ӳ�l\ Ө��BI;�p�A��7��:i#]W�*t���?�,�����K�ſ'���䫉Fm�7'g��l?'�v���\�"v@�j[mUC��[��ITk�C���^V
�-�U��3C܇����(pTB��/U�}lI��Ah��E��v#U���:��ο&)�T�A����-X���C=e��G�k(�d��������#�dHc>��w�"�LCg�3K�jnD|)�rp��Gq����w�>.�sT�ߥ�h�<t<N�g���f����+�u��SmF�2�P>�J�Y���ƈ��B7���K R�5Q��B���UG���<�&��~��`3�^�;4���02Uƿ�y��H|�����U���Ov����k�&��H��/y��&ˬL.�K8��H��r�V��g���GU��qrAՏ�ne�5���P]��|�=� ����B
�H����OT���&��Ö�i��4Oq=P9w���E��VTf��k{K��Y�)}�穚������qWq��E�i"	�g���:��k���iϹ��XH{F�I�_���3;G\'��ZJ˙�`��n�5��E�NԨ8Л-]G�%��p6�L�ʒq��W<��{科{Ç��@]�����X�PxvD4�Ue3���o�R@�+�/�����ܑ�3{?<��'w����j���f�R i�	0����Մ�%�:i;���pC��W�PKz$+ K�I3�%�qVnO��ǫۡg=�׉O�͂�d%�HU����塪A��;K��\�ޟv1�i�gΣW���s;E�`�@y�W�p@����!��4b�l�o�G��.Gw
#XE`��Q�p�&����.T�x�:�޺����٩���H���6�s�z���R��@����D�
��9���+D�>2�6�dm�Cc�G~�n,0�>uٔ�U�F@	ʝD;�f�)�adY(�f��_-��諣P�8}s2i@�D�[X��2NP��ע��U趣���(�QB�$m�`�gq&��x�{���{��z�	��=�^4�
#���Қ1`z�US��J�H)�.v>�n`��[�y�W��w�p/f>�QP�"�%n�y�v� qp��I���ƼWܿ���wOSú�R?3|�5��Fg:VM{�BK`��>���~h�k>�%�=���HD��g��)x��TA�]ڟ/��Ҝ�U�^˜�W��W�����8�w��a�B�Tږӵ�b�;�����kD[ONc_����>��Ƣa)�J����f�mS=T �Gំ��(�)r��&"�����x���xd)xf�� Ҋ�$!5(���_���E�S`�&���穣���:#������uX���&������T�p�ɤ7��P*��B=7=²�fd���.�s�P��c~��Y̗ �v{�p�g�lI�_�Iδ�S��F��s�gE�3{.�T/AC'GYJ w����	�9�S��foS�7��l��B�o� �������C�/�S+�IC��%'�=C�>Y��ld�{��+��GbN�[ �� �$g��+Q4�~4�W��8Od�\���!e�SSF>(�ך>A>���9��K�)���K����<�V"��+��S{
wE�+�/�cnh@�������TBD>5k��GJ���eщ�� �%�.������0�^�f`��}w(�"�y'p3�vF�녦�@ր��f뗩p��U吥��3�R�T���V�FFzDꎐH�:�<�<�h�R)�ۗ'|d�O��{2p����$���^�� v4P�MBqnZ�&��b:�E��خ�G�V;c���f( �3�}|d�_	g�����1W�m�W)N��2�ߧ�b"������B�9 "7	�5��M-5F(���vuk��T(�8r6��6K|ʕ��c�!�,{M�7���M�X���5O%ȝw7O��k�O��ن�o���e�`�)�@�}+&��k�"���e�1Ii)����{ڣ�����\�s]��$0#��ui?��khV���<�=k�to�5��5L����
��k�w��Ne��CC�"�ێ~x�0C�q���\�B,뙖��)B��M�lO���*�%�����ͪ��MV���tԥ��}���3��P�и�⏥��}�b̺�-��j�V��pI����6�9�?�_[J��5M �A/�9��A�8�ϫ��Ŋ�C*�c����G�SY�X����Ґ, ���L�ӡ�먮��vx�V���).�c=�!��3��8�R�oq�̔&B1�/KS���. [��=�u�b�1��I!�E���?�V7B��B����[,m��n��zZ�>9�>���S�A�ܮ�����=�l��k�1}#��>�NC=>v��f��Z�e�j��n!{?#W��9ؒ��r�X���=kv���� �b�nH� ����PXY������)cc�������d���W �=�g9��������1��*^{"���po�#�ۑ'�b�	����	����î�p�I�Y�#,]�jCG7b!��oܴ�L�Ն�����;�X�I�¤��^A����i~�q� ����Ŵ�u��~�8nJٟ�����=��N��\�G�����i9��Z�sVO�)���$�3����*L~9�x.�[Ky��|�ѝ������,�j*]��M����?�i0򥏐|�װTc�cm^�&+�a�_��$�
A!�W����a����\h� ��.���X������A�����
��G4��ͻ�.��H�+k�ܟx�VkJK♬�����تa2��քl�3�O�3.�"˼#�ު�W� +^�B̀��*:��O��l��SX��>B��t������=�^��-̜F3��?�A��އm�GJ��
'�tBD!�1N���^�]��#T�	��oC���":�e��1�(bR)���l�§���'È��@!/��m#�<�R����hAO�G�%��#��+����K*���A�F���r���)�#��+�Q&B������9�]�#t��㕒�t�N�N�Q��V�u�����P�	�/��\v��JA ^�Nz=�*ZȔ���Fp9>͈�R�*z�I�#�j9P	W����� ��e�+�_�q^K�ٺB�o�Ê`0=���r!JiT��qg�"��Ng�#u��� ��=�m��u� � W����\A.ԐG���g-f7}tI�m-؜*^����y���|�Г�x��2Z��:��P.���l��턩�oDK���<~$ddaK���h�M�&�{H�F7Y�
������h<�`ӽ�g�&�Zl���&�?����m�id;#���n楉�N�M�f&[l��~���9��V5���#�W:�4�v��hP�����v�j��\�-�>�a�f9�W䙫h�LL&ԝO*V#��F @��u��n�V���%�Ut~����zz#`9�(��M�q�\����G�t��*����w����-/2Rn���,�[�6�U����q+Q�'�*A�Iy �oqH�g�s]R�ԁ`�k)��*�tr���G���H;�b�X�������ɼYl&2)�L��!��yBco���k)+�����k-F��a�Z�{`Tg�wL�
0!��K}�F���U(XJ�� 4|�Ia�����d�Uc�����h�v���n�!�~��6�e�O#��:�Ϧθ/���\	�B��j�K��bj}�j�������QA)�i�?�%����=DLr�̞4"��@+�%n����mN��¾�D��L�"������%�¿�����وF=�]� q�bN���Y�,*5u��i�Z�a�?�2j}9�����l�t��s_�����Nc���oM��2���A�Z�(b� ��� �?q�ۉ�M2�1�J�v�k[��.�+p����	Ɇr�<>TR�̇,��6�	������P⯵W\�1@��<B>�L�G��l\�p�E�]
��@�@Ɯ��WBj�v;�k�,�?5|���255a��% ���*ۿ�j;@���	��`(â:S%��a�����$h�b��������6x��#= 5�NvH�@a�"h��L~R�mv	��+N��ޠ�ȁ�;8S���4㫢��j%ƀ�u����5�Z%��ڢ�����r(��0 0���J���6���?ȻOGe�KHHr�Qp���YG��#�D�����m����HJ"��6Й�$�K����K���Z/'/�ƭ�q�]g��De'F|���r���zug5ͥ9���C����g�i���|�j�h8�n=by�!�r�{����C��35D�r�����j�H��MOm}h�9�y_����R�����M��2���J+5�"�l�/�?f��o�Uj_���2�l؊ƣ�zm;��Q�Tު��´��~Z�(�y��r�-��Avg�Z�c� )i]��83��cE����hE��vo�^������4�p�O��=
�q��.��%\d/��C?��(1A=Hr�P;׻��۩k�q��g�r�0�@��(|�`#��|�I���W��ߔn"���f.Gf��>�f<������>����vqN�;����FK@h�cw�o�9Q�<�JN_�&1V �Z��P��_��'�]�h����U��6��e���4�i?�Qs�6p��r"����h�,��X�b��*.�n�I��m��rr6���6��=Gv��V�Z{P�Ԑ:A ;�Z����S5-~��t�y�>�I(L�)�Y��6Ji��.��2Z�z"L��&.,C!������Pwx��&�}\.���9���"�X�g�R��"���jG\�+7����6��)�H��J����y�u �Cke梉G�k[��X'n�Qi�q(��7���37�A�p��gUH��(�䜤  ��m�U�cNK&A�OwB�!�7_��܀c5¿�(�(�+�Ut��O���3��0z��ɌN��?X|R���2p�A�E��ºz�L�X��￸w�G��L@�\z�)�(�鿡�`�J�<O�7�9j�4Dm<jO�u<O�a%�׬�h�x�Z9�3��:���V��^E<���S��V�(�������e���(ߟ�9G��;�7�����Е¼l�/RiY��/$w�D���H.Lc��uQ�� yuK�����KP`��E���E;T�Hg)fչ^�כ�jTo	���WG�m��ȸ�5-���~��M�V���l<�6��N�"	
�gZ��3FO�q3;4ץ�٘KjѠ��(}���N��Y��i]D$DM�!Ι�!a苝E�ԫ����Y�Pk� �h���׆�~�ј1�Q�����F� �\����+�v�Y9i�tҧ��O,������~���rMR?��o��mIc|�Bu�OţFJ��r�ћj�Rd�Ȕ�|�5E>�媒��4z�s�!�J{}{^C�f9"]p�<R�ӎ��� �'��q�[�~�9��, ����1S�|�}%@�jbN&��)J�J�J�tl7$�*M�
�B�.�<�^�e+@���������i�9��cH��֒�	쒒b�L{��~���Y��=�j"%�b0N�̝M�du���d�*��2�����@/�l[@6H/�G]�y��A��)���UZ'�n��U7�����	&"��`�Y2%���S'�����aa��������Ba�́P�� 6ڹ����ztJ����[�j!�VE�=B?�\��G�0ǟ!�^�PVw�w6/6�+�����GM���I���v Gѧ�L����b��X���9jt��9$Љ������<���kѽ�"P��N�m6����v����p����;u��D/�@��ة�8�G�����|�҉���� �x7��jN&e|E1�o��X懑.2g��w�	(B]!���@���%sQw�F��O���r�Dw#7"͈�;%����v팜I������@X<_11�ِ�au�	����੊��$��.,�ƙ�W��������`_}13+0�a���tu�̭/��������q0(���ƌP�1[��v�/�zW`��e3�ՇK��/�����M�����؇��NX���5cW2l�T����;?c�q�p}|���9��¥*�,���0a�p��鯣��)P.��C.�k��Е���)�r*��³�{�ߕ����+*��pL�=e���G	�K�����bƨ+vSp����H��V�M �i���2l��1H�RV� Ռ� �;�>!h1gg�����&$?J)��6zW<�CBP�|�@����]�з޿w����ڛ+-'�g�4;q��.qh����oTI� R�tɔGI������暘?L"��92����.f�[Z���mP�ܲ��uw�V��R��j	'J֪��[<O@�܉��}�SW��{ �o]p;�����
ŕA=P��:E��&׊m\�y���: �9�ܸ�#�#������$�v�"�mVR�D|0IG��j������G
9G�\�8�������`�	nU����3Z��S`8��U��}C�X:���h���T>n������:��,%R�F���h��sG�[Fq��F{�>�K�J�L��
b�V>��K�@�.������j�����M	��טm�6��d�3�ѯ�|^�E46^ue�I�(��$������}&�}E�.��mo;w��X�:�Wg�	�͉]O�˭*�Z�|�m���YiAz��A�=cw��ɫ<�I|(U]4&�@�*׿W�������Ȫ|b���;���<�]b̶-P�I�Xg-��5b��9_������8hPq���Ø9��*ST0�+rڌ�J+{�ѫd)MU�*��go:9B<��8p��vJ�7+!]��ڛj�Fߣw ���s����U{����u��q-p���/��.�g#��W���*4w�e�_�V}�xs��t?�P@P)\��|�Q>�˃(�6|={���鰃߉*��u�dl��;U� ��l��	�\�������y��u��A��^A~���Z��:����Cab�y���ڽV���T���rh�Ó������rI���M&L��au-F,�l�O�j�.�?���5�6c�ۈ���S�:���{u���r�.�z��h�.�g�L���;Q%#��N�}�$��� �����֚M��&~�Z̛��=�MoJ�M|k��$����&�9*�<���6퓫���]�-U]��x�;h�S,3��r~\�E
��$�7�f�8�(2O�3\�S�,���(��%J�^����ߪe�fى��%��p�r��2�g��S_��h3"lh���G(0�?�F/����(�.�J`6'����5ԅ�ѕ��V����\}��^\,��h��H>�㷩|����(β���F���Q���IhDrR8��(�_�z��g2T�#za<��H���޳O��fb�ә�@�吿��u�d!�b�u��P=2��,V�6���h�TZcS�g��;Z����ōݜ  ���Em%z@��iu�hV�*z��^Еc�#�2K��O�f�i�Fd��m�h�k�#�zd���Y{[�Q��y�r�hzc��0��&��'.��� ΂A�9���c���(��S�˚j�;}g�H�6ڥj�`U�z�@~_+��qC����Ŋ|�Z�wj^zI����ˢ��#hd Hi�ظK Mn�9|^�m�GL��c�]��	���a-�O��	�E��\�c׻WFe��R���.()�FL�q��a����`u�1����/�9���_������f��Ю�_uҶW���Q��9n暢�r�R�2S���OL��'hT�t���-ΠaN�HTsB��.j$��Ϫy���(�����q5XҼ&'l�|A�&b��y�ߖ�f%�>�`���?>���ow�oQȾ���-�8飽l� �2NղB��+[�[j��P�1��+��W�V7u�}�|�!R�G���3�x�\MP;Ld~������j Ot�@���Eu�3�A-�Z4�5CY攃�vy��X�(�+I�����Kw�p���}?jӣ������� }E��J��a���x4Z�>��E�'t�z�̿D/_-�\nm��-��c����bVi0o��e-=�y�ѕc-�r8ۨ�iFc��˿�N���1��������x�����uC��O�4���o��l�"Cr��@�b,�,:���f��]8T���]:�pc����2��Jѓ񎐑���o��Di#�M�Ȇ9�`�T��)h��-h��ړ+��}w� 
��)1^>�K�dz��
�G/a�5mU�&A�5뉊!^Q��`o������jN�Kض�HL"�	$v���(��,8�TA���]������*�>�+���Z̘��(�7r�C6ņ^�e�%p;��k�̸��Nrց&0��T��Tr@��{��֟�?����O'p�D�p��c[��qV����f�<*G��u9���I�t^>P��'ݰ��~���p��3*���X� ��!�n���Г�?%[t����CZǏ�e~'��dB��9� �h��'9�J�����0��ֲdZaNٔS
SV�:�=7}.�D6�bԖ
 �Q��`��;dz�e�{!�{6E[+�v�����jͳ&�oNd7!�@��B2;�D��P����E/���(0��G�$���~"]b f�6�MM�c
��׾q.�t���޴�̳ĞR;B����r������E�x�}"���A�)�%�@�ڀ#�E'�{�M������� V��l�ccl�Nc~#sj߄��g�=�9��]��\"����_4t��J+�'����G���-�k��^%J�5�n���d!�7�Gd�ha��-������sq�q��E�R��T�Zu�~��:}Qv����c`����*�^cNJ.`x���B����vz�q!M�2���[#�T;� r	��"��u����"0���_� C�ñ��1�+�>O�&��N)2�B��y��ھ^<���lTti� �� Z��?���w\���+Ɛ�3�"-]��yղeS�c���|�>g8�Z=���6u�M���f��7pPT�g�[+%��cb���sR������*U�^���P"P:��>b4H������1]Zq�̷�yT�t �s�d���.���1�
�ͮa��S�!v��!vAL��2�h��4<�`�HL�w�&���@� �	�������	z��D%�ם�#�Z;�@̔g.�˖3\��@�X�0zs���'C��q�� �������Y��������R�)F}B���Y���|���	'"����� �4��\�:����%:G�����5��ĸ���o�*9�r�S�ʕ�G"b0ʨ����K���.�.��Y��[OF�^dN���6�PF;K	����`[p����TpA�џՑ�P�+q�S%w�_{^�^(�)�SN�mN�i�����!,e��2��Y�!H>����������H.���"PE��?u��		9�{��/��9o�%9����*$#��F���|��!OSޞ٢��B��n`'��6d�$L�g���f��(]q��vۮ����:�]z�fb�pR�:��������7��r�GÓ!|�ZǤ��#�M��|�&�'ys#����+"���	�W����ɟc���}�Q�@Ls�D1���z*�b{q��%:eY� ��zU��Qb�I�h m� ��H��s.�z����V+Dv�΢��ʿC��4?oAs�@q�t�O�����ᄄ'Z9�� j�Ϟ�/k��o���,Bg�����v�+5�`����Q(m�z�m�B�����1]O[}[�4��Y�-��0�����W�P����L|?&�Bc���"�Tͳ������a�:W�@;@HI<��E�k����r#���}�],#��MD<�B��P�ac����Y���GTy��U�Qy6B�u�B�n�����Kd<|ݫb
�&�3q<���\��ڲ����~*���4��M�ui9��M*���b[S$YV���8�O�*p��O7��WDv>ץ��z�Gr��~�\nY\��7����}���8��p��l���}8~�]�(�9eLqu�t�g����^XC������Q�"hH�a&�ɟ0��6���Tl
m��9�������>P��֊M�$B�&ũ��*�b�)���T%s�)�6I{_k�R�d�O�-�Ź���T��W�	���N�鑶����[K���a!���'5�ep@PF�,��h�D�'��d����ȱ��z�OO/����`I�Ӗ�[���1;m%�Vך!i�f���Kff3�}�B�z���T΍�%jy���F�G+�C�r[�>P�����;��J�@��\#�a�����E�z��)�R��m��A�9���"�c�k�z��A�5��V5�m�P���)�����m=��z`�Km%�*`��(h��B�Xg%�=�ӀUߥ�Hlb�lr���n}^=t7v��ڮ��ؕցx��ZO�������PB��W��$����oN��ԩn^Q��vO�H�D�B5���&��L�_��6�1���O�07k_�ǿ��`���r���]�W֥���Z����Ns��K����	�k}V�!j�������S�x����/�8T#�v�S�����ܢD�~�KL�� �r�!�EY�J]�����b����;5�g��� ^t�&⟜Mx �OЄi[!7�q*��t��ZN�|*��2^�U=-�@{�"���⺞N����N�@#~�[=L&$�IԘ�,X3BB��A�Zk�eo�C�sT���G^J�v�Ӷ��E�;3�g�vHF[�q�����zu�~�K���f��۰[���E��%6w�e���P�D��Wo��}���)f@~���#,4.�����E.���pi�^�.��lG�%s+��u����.`�]s�U�#�3��̥�.�ю+o^Kׂ�0��P�������ҧg���ɱ�O��5f�@� J�W����^hט�UX|�dWK�u9n<��"�w�L_��*��h����*��^iw��� �,���ɽ�>��P�#�Fo�D4����m���"�x��E>�#�}r�Lb�{~���[�k>P[�09I��:��u���� �E=Tpq�,�:��i�l>3	� �|�(������8V�ogfT�Ȗ���ײ���N�k�$��k�<d�?1n���3!���껉R7����/���8jvE4Q�=�e:�;A�� ���[�6��&+�ޕ�U~��x���mL%��Ua=�^z�^������sNR4�;���+-�n��r���@a�=�:�kR��ǐf}\���Q0�y D� �aSd�\��eo�AY�SI�@RB,��PBb_��W��R����o!�5��27*�x�z$��8���|O����� h�;4���eRϗ��8�A>�}�V��	b��D}g�I$�O �Xx49�,#ܱ�i��r���t�6���ǉ-R6�-ğ��B8<���ߍ�'E�\�v�(��9Ҥ>�� ���u��w��t����h�6�%�K��j��Z�5+�?�yƟ5�b�H��k$�-��z�]I�d��s�\ �ܒ���T��E��k6ܮ�^˳���E�v�p2H�u7sÊ�X�;��댠S{�L